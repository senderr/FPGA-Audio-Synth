module sine_wave_generator (
                            clk,
                            enable,
                            fn_in,
                            signed_bit,
                            out
                          );

  input clk;
  input enable;
  input [10:0] fn_in;
  input signed_bit;
  reg [31:0] sin;
  output reg signed [31:0] out;

  always @(posedge clk) begin
    if (!enable) begin sin <= 32'b0; out <= 32'b0; end
    else begin
      case(fn_in)
        11'h0: sin <= 32'h00000;
        11'h1: sin <= 32'h000032;
        11'h2: sin <= 32'h000064;
        11'h3: sin <= 32'h000096;
        11'h4: sin <= 32'h0000c9;
        11'h5: sin <= 32'h0000fb;
        11'h6: sin <= 32'h000012d;
        11'h7: sin <= 32'h0000160;
        11'h8: sin <= 32'h0000192;
        11'h9: sin <= 32'h00001c4;
        11'ha: sin <= 32'h00001f6;
        11'hb: sin <= 32'h0000229;
        11'hc: sin <= 32'h000025b;
        11'hd: sin <= 32'h000028d;
        11'he: sin <= 32'h00002c0;
        11'hf: sin <= 32'h00002f2;
        11'h10: sin <= 32'h0000324;
        11'h11: sin <= 32'h0000356;
        11'h12: sin <= 32'h0000389;
        11'h13: sin <= 32'h00003bb;
        11'h14: sin <= 32'h00003ed;
        11'h15: sin <= 32'h0000420;
        11'h16: sin <= 32'h0000452;
        11'h17: sin <= 32'h0000484;
        11'h18: sin <= 32'h00004b6;
        11'h19: sin <= 32'h00004e9;
        11'h1a: sin <= 32'h000051b;
        11'h1b: sin <= 32'h000054d;
        11'h1c: sin <= 32'h000057f;
        11'h1d: sin <= 32'h00005b2;
        11'h1e: sin <= 32'h00005e4;
        11'h1f: sin <= 32'h0000616;
        11'h20: sin <= 32'h0000649;
        11'h21: sin <= 32'h000067b;
        11'h22: sin <= 32'h00006ad;
        11'h23: sin <= 32'h00006df;
        11'h24: sin <= 32'h0000712;
        11'h25: sin <= 32'h0000744;
        11'h26: sin <= 32'h0000776;
        11'h27: sin <= 32'h00007a8;
        11'h28: sin <= 32'h00007db;
        11'h29: sin <= 32'h000080d;
        11'h2a: sin <= 32'h000083f;
        11'h2b: sin <= 32'h0000872;
        11'h2c: sin <= 32'h00008a4;
        11'h2d: sin <= 32'h00008d6;
        11'h2e: sin <= 32'h0000908;
        11'h2f: sin <= 32'h000093b;
        11'h30: sin <= 32'h000096d;
        11'h31: sin <= 32'h000099f;
        11'h32: sin <= 32'h00009d1;
        11'h33: sin <= 32'h0000a04;
        11'h34: sin <= 32'h0000a36;
        11'h35: sin <= 32'h0000a68;
        11'h36: sin <= 32'h0000a9a;
        11'h37: sin <= 32'h0000acd;
        11'h38: sin <= 32'h0000aff;
        11'h39: sin <= 32'h0000b31;
        11'h3a: sin <= 32'h0000b63;
        11'h3b: sin <= 32'h0000b96;
        11'h3c: sin <= 32'h0000bc8;
        11'h3d: sin <= 32'h0000bfa;
        11'h3e: sin <= 32'h0000c2c;
        11'h3f: sin <= 32'h0000c5e;
        11'h40: sin <= 32'h0000c91;
        11'h41: sin <= 32'h0000cc3;
        11'h42: sin <= 32'h0000cf5;
        11'h43: sin <= 32'h0000d27;
        11'h44: sin <= 32'h0000d5a;
        11'h45: sin <= 32'h0000d8c;
        11'h46: sin <= 32'h0000dbe;
        11'h47: sin <= 32'h0000df0;
        11'h48: sin <= 32'h0000e22;
        11'h49: sin <= 32'h0000e55;
        11'h4a: sin <= 32'h0000e87;
        11'h4b: sin <= 32'h0000eb9;
        11'h4c: sin <= 32'h0000eeb;
        11'h4d: sin <= 32'h0000f1e;
        11'h4e: sin <= 32'h0000f50;
        11'h4f: sin <= 32'h0000f82;
        11'h50: sin <= 32'h0000fb4;
        11'h51: sin <= 32'h0000fe6;
        11'h52: sin <= 32'h00001018;
        11'h53: sin <= 32'h0000104b;
        11'h54: sin <= 32'h0000107d;
        11'h55: sin <= 32'h000010af;
        11'h56: sin <= 32'h000010e1;
        11'h57: sin <= 32'h00001113;
        11'h58: sin <= 32'h00001146;
        11'h59: sin <= 32'h00001178;
        11'h5a: sin <= 32'h000011aa;
        11'h5b: sin <= 32'h000011dc;
        11'h5c: sin <= 32'h0000120e;
        11'h5d: sin <= 32'h00001240;
        11'h5e: sin <= 32'h00001273;
        11'h5f: sin <= 32'h000012a5;
        11'h60: sin <= 32'h000012d7;
        11'h61: sin <= 32'h00001309;
        11'h62: sin <= 32'h0000133b;
        11'h63: sin <= 32'h0000136d;
        11'h64: sin <= 32'h0000139f;
        11'h65: sin <= 32'h000013d2;
        11'h66: sin <= 32'h00001404;
        11'h67: sin <= 32'h00001436;
        11'h68: sin <= 32'h00001468;
        11'h69: sin <= 32'h0000149a;
        11'h6a: sin <= 32'h000014cc;
        11'h6b: sin <= 32'h000014fe;
        11'h6c: sin <= 32'h00001531;
        11'h6d: sin <= 32'h00001563;
        11'h6e: sin <= 32'h00001595;
        11'h6f: sin <= 32'h000015c7;
        11'h70: sin <= 32'h000015f9;
        11'h71: sin <= 32'h0000162b;
        11'h72: sin <= 32'h0000165d;
        11'h73: sin <= 32'h0000168f;
        11'h74: sin <= 32'h000016c1;
        11'h75: sin <= 32'h000016f3;
        11'h76: sin <= 32'h00001726;
        11'h77: sin <= 32'h00001758;
        11'h78: sin <= 32'h0000178a;
        11'h79: sin <= 32'h000017bc;
        11'h7a: sin <= 32'h000017ee;
        11'h7b: sin <= 32'h00001820;
        11'h7c: sin <= 32'h00001852;
        11'h7d: sin <= 32'h00001884;
        11'h7e: sin <= 32'h000018b6;
        11'h7f: sin <= 32'h000018e8;
        11'h80: sin <= 32'h0000191a;
        11'h81: sin <= 32'h0000194c;
        11'h82: sin <= 32'h0000197e;
        11'h83: sin <= 32'h000019b0;
        11'h84: sin <= 32'h000019e2;
        11'h85: sin <= 32'h00001a14;
        11'h86: sin <= 32'h00001a46;
        11'h87: sin <= 32'h00001a78;
        11'h88: sin <= 32'h00001aaa;
        11'h89: sin <= 32'h00001adc;
        11'h8a: sin <= 32'h00001b0e;
        11'h8b: sin <= 32'h00001b40;
        11'h8c: sin <= 32'h00001b72;
        11'h8d: sin <= 32'h00001ba4;
        11'h8e: sin <= 32'h00001bd6;
        11'h8f: sin <= 32'h00001c08;
        11'h90: sin <= 32'h00001c3a;
        11'h91: sin <= 32'h00001c6c;
        11'h92: sin <= 32'h00001c9e;
        11'h93: sin <= 32'h00001cd0;
        11'h94: sin <= 32'h00001d02;
        11'h95: sin <= 32'h00001d34;
        11'h96: sin <= 32'h00001d66;
        11'h97: sin <= 32'h00001d98;
        11'h98: sin <= 32'h00001dca;
        11'h99: sin <= 32'h00001dfc;
        11'h9a: sin <= 32'h00001e2e;
        11'h9b: sin <= 32'h00001e60;
        11'h9c: sin <= 32'h00001e92;
        11'h9d: sin <= 32'h00001ec4;
        11'h9e: sin <= 32'h00001ef6;
        11'h9f: sin <= 32'h00001f28;
        11'ha0: sin <= 32'h00001f5a;
        11'ha1: sin <= 32'h00001f8b;
        11'ha2: sin <= 32'h00001fbd;
        11'ha3: sin <= 32'h00001fef;
        11'ha4: sin <= 32'h00002021;
        11'ha5: sin <= 32'h00002053;
        11'ha6: sin <= 32'h00002085;
        11'ha7: sin <= 32'h000020b7;
        11'ha8: sin <= 32'h000020e9;
        11'ha9: sin <= 32'h0000211b;
        11'haa: sin <= 32'h0000214c;
        11'hab: sin <= 32'h0000217e;
        11'hac: sin <= 32'h000021b0;
        11'had: sin <= 32'h000021e2;
        11'hae: sin <= 32'h00002214;
        11'haf: sin <= 32'h00002246;
        11'hb0: sin <= 32'h00002278;
        11'hb1: sin <= 32'h000022a9;
        11'hb2: sin <= 32'h000022db;
        11'hb3: sin <= 32'h0000230d;
        11'hb4: sin <= 32'h0000233f;
        11'hb5: sin <= 32'h00002371;
        11'hb6: sin <= 32'h000023a2;
        11'hb7: sin <= 32'h000023d4;
        11'hb8: sin <= 32'h00002406;
        11'hb9: sin <= 32'h00002438;
        11'hba: sin <= 32'h0000246a;
        11'hbb: sin <= 32'h0000249b;
        11'hbc: sin <= 32'h000024cd;
        11'hbd: sin <= 32'h000024ff;
        11'hbe: sin <= 32'h00002531;
        11'hbf: sin <= 32'h00002562;
        11'hc0: sin <= 32'h00002594;
        11'hc1: sin <= 32'h000025c6;
        11'hc2: sin <= 32'h000025f8;
        11'hc3: sin <= 32'h00002629;
        11'hc4: sin <= 32'h0000265b;
        11'hc5: sin <= 32'h0000268d;
        11'hc6: sin <= 32'h000026be;
        11'hc7: sin <= 32'h000026f0;
        11'hc8: sin <= 32'h00002722;
        11'hc9: sin <= 32'h00002754;
        11'hca: sin <= 32'h00002785;
        11'hcb: sin <= 32'h000027b7;
        11'hcc: sin <= 32'h000027e9;
        11'hcd: sin <= 32'h0000281a;
        11'hce: sin <= 32'h0000284c;
        11'hcf: sin <= 32'h0000287e;
        11'hd0: sin <= 32'h000028af;
        11'hd1: sin <= 32'h000028e1;
        11'hd2: sin <= 32'h00002913;
        11'hd3: sin <= 32'h00002944;
        11'hd4: sin <= 32'h00002976;
        11'hd5: sin <= 32'h000029a7;
        11'hd6: sin <= 32'h000029d9;
        11'hd7: sin <= 32'h00002a0b;
        11'hd8: sin <= 32'h00002a3c;
        11'hd9: sin <= 32'h00002a6e;
        11'hda: sin <= 32'h00002a9f;
        11'hdb: sin <= 32'h00002ad1;
        11'hdc: sin <= 32'h00002b03;
        11'hdd: sin <= 32'h00002b34;
        11'hde: sin <= 32'h00002b66;
        11'hdf: sin <= 32'h00002b97;
        11'he0: sin <= 32'h00002bc9;
        11'he1: sin <= 32'h00002bfa;
        11'he2: sin <= 32'h00002c2c;
        11'he3: sin <= 32'h00002c5e;
        11'he4: sin <= 32'h00002c8f;
        11'he5: sin <= 32'h00002cc1;
        11'he6: sin <= 32'h00002cf2;
        11'he7: sin <= 32'h00002d24;
        11'he8: sin <= 32'h00002d55;
        11'he9: sin <= 32'h00002d87;
        11'hea: sin <= 32'h00002db8;
        11'heb: sin <= 32'h00002dea;
        11'hec: sin <= 32'h00002e1b;
        11'hed: sin <= 32'h00002e4c;
        11'hee: sin <= 32'h00002e7e;
        11'hef: sin <= 32'h00002eaf;
        11'hf0: sin <= 32'h00002ee1;
        11'hf1: sin <= 32'h00002f12;
        11'hf2: sin <= 32'h00002f44;
        11'hf3: sin <= 32'h00002f75;
        11'hf4: sin <= 32'h00002fa6;
        11'hf5: sin <= 32'h00002fd8;
        11'hf6: sin <= 32'h00003009;
        11'hf7: sin <= 32'h0000303b;
        11'hf8: sin <= 32'h0000306c;
        11'hf9: sin <= 32'h0000309d;
        11'hfa: sin <= 32'h000030cf;
        11'hfb: sin <= 32'h00003100;
        11'hfc: sin <= 32'h00003132;
        11'hfd: sin <= 32'h00003163;
        11'hfe: sin <= 32'h00003194;
        11'hff: sin <= 32'h000031c6;
        11'h100: sin <= 32'h000031f7;
        11'h101: sin <= 32'h00003228;
        11'h102: sin <= 32'h0000325a;
        11'h103: sin <= 32'h0000328b;
        11'h104: sin <= 32'h000032bc;
        11'h105: sin <= 32'h000032ed;
        11'h106: sin <= 32'h0000331f;
        11'h107: sin <= 32'h00003350;
        11'h108: sin <= 32'h00003381;
        11'h109: sin <= 32'h000033b2;
        11'h10a: sin <= 32'h000033e4;
        11'h10b: sin <= 32'h00003415;
        11'h10c: sin <= 32'h00003446;
        11'h10d: sin <= 32'h00003477;
        11'h10e: sin <= 32'h000034a9;
        11'h10f: sin <= 32'h000034da;
        11'h110: sin <= 32'h0000350b;
        11'h111: sin <= 32'h0000353c;
        11'h112: sin <= 32'h0000356d;
        11'h113: sin <= 32'h0000359f;
        11'h114: sin <= 32'h000035d0;
        11'h115: sin <= 32'h00003601;
        11'h116: sin <= 32'h00003632;
        11'h117: sin <= 32'h00003663;
        11'h118: sin <= 32'h00003694;
        11'h119: sin <= 32'h000036c6;
        11'h11a: sin <= 32'h000036f7;
        11'h11b: sin <= 32'h00003728;
        11'h11c: sin <= 32'h00003759;
        11'h11d: sin <= 32'h0000378a;
        11'h11e: sin <= 32'h000037bb;
        11'h11f: sin <= 32'h000037ec;
        11'h120: sin <= 32'h0000381d;
        11'h121: sin <= 32'h0000384e;
        11'h122: sin <= 32'h0000387f;
        11'h123: sin <= 32'h000038b0;
        11'h124: sin <= 32'h000038e1;
        11'h125: sin <= 32'h00003912;
        11'h126: sin <= 32'h00003943;
        11'h127: sin <= 32'h00003974;
        11'h128: sin <= 32'h000039a5;
        11'h129: sin <= 32'h000039d6;
        11'h12a: sin <= 32'h00003a07;
        11'h12b: sin <= 32'h00003a38;
        11'h12c: sin <= 32'h00003a69;
        11'h12d: sin <= 32'h00003a9a;
        11'h12e: sin <= 32'h00003acb;
        11'h12f: sin <= 32'h00003afc;
        11'h130: sin <= 32'h00003b2d;
        11'h131: sin <= 32'h00003b5e;
        11'h132: sin <= 32'h00003b8f;
        11'h133: sin <= 32'h00003bc0;
        11'h134: sin <= 32'h00003bf1;
        11'h135: sin <= 32'h00003c22;
        11'h136: sin <= 32'h00003c53;
        11'h137: sin <= 32'h00003c83;
        11'h138: sin <= 32'h00003cb4;
        11'h139: sin <= 32'h00003ce5;
        11'h13a: sin <= 32'h00003d16;
        11'h13b: sin <= 32'h00003d47;
        11'h13c: sin <= 32'h00003d78;
        11'h13d: sin <= 32'h00003da8;
        11'h13e: sin <= 32'h00003dd9;
        11'h13f: sin <= 32'h00003e0a;
        11'h140: sin <= 32'h00003e3b;
        11'h141: sin <= 32'h00003e6c;
        11'h142: sin <= 32'h00003e9c;
        11'h143: sin <= 32'h00003ecd;
        11'h144: sin <= 32'h00003efe;
        11'h145: sin <= 32'h00003f2f;
        11'h146: sin <= 32'h00003f5f;
        11'h147: sin <= 32'h00003f90;
        11'h148: sin <= 32'h00003fc1;
        11'h149: sin <= 32'h00003ff1;
        11'h14a: sin <= 32'h00004022;
        11'h14b: sin <= 32'h00004053;
        11'h14c: sin <= 32'h00004083;
        11'h14d: sin <= 32'h000040b4;
        11'h14e: sin <= 32'h000040e5;
        11'h14f: sin <= 32'h00004115;
        11'h150: sin <= 32'h00004146;
        11'h151: sin <= 32'h00004177;
        11'h152: sin <= 32'h000041a7;
        11'h153: sin <= 32'h000041d8;
        11'h154: sin <= 32'h00004208;
        11'h155: sin <= 32'h00004239;
        11'h156: sin <= 32'h0000426a;
        11'h157: sin <= 32'h0000429a;
        11'h158: sin <= 32'h000042cb;
        11'h159: sin <= 32'h000042fb;
        11'h15a: sin <= 32'h0000432c;
        11'h15b: sin <= 32'h0000435c;
        11'h15c: sin <= 32'h0000438d;
        11'h15d: sin <= 32'h000043bd;
        11'h15e: sin <= 32'h000043ee;
        11'h15f: sin <= 32'h0000441e;
        11'h160: sin <= 32'h0000444f;
        11'h161: sin <= 32'h0000447f;
        11'h162: sin <= 32'h000044b0;
        11'h163: sin <= 32'h000044e0;
        11'h164: sin <= 32'h00004511;
        11'h165: sin <= 32'h00004541;
        11'h166: sin <= 32'h00004571;
        11'h167: sin <= 32'h000045a2;
        11'h168: sin <= 32'h000045d2;
        11'h169: sin <= 32'h00004603;
        11'h16a: sin <= 32'h00004633;
        11'h16b: sin <= 32'h00004663;
        11'h16c: sin <= 32'h00004694;
        11'h16d: sin <= 32'h000046c4;
        11'h16e: sin <= 32'h000046f4;
        11'h16f: sin <= 32'h00004725;
        11'h170: sin <= 32'h00004755;
        11'h171: sin <= 32'h00004785;
        11'h172: sin <= 32'h000047b5;
        11'h173: sin <= 32'h000047e6;
        11'h174: sin <= 32'h00004816;
        11'h175: sin <= 32'h00004846;
        11'h176: sin <= 32'h00004876;
        11'h177: sin <= 32'h000048a7;
        11'h178: sin <= 32'h000048d7;
        11'h179: sin <= 32'h00004907;
        11'h17a: sin <= 32'h00004937;
        11'h17b: sin <= 32'h00004968;
        11'h17c: sin <= 32'h00004998;
        11'h17d: sin <= 32'h000049c8;
        11'h17e: sin <= 32'h000049f8;
        11'h17f: sin <= 32'h00004a28;
        11'h180: sin <= 32'h00004a58;
        11'h181: sin <= 32'h00004a88;
        11'h182: sin <= 32'h00004ab8;
        11'h183: sin <= 32'h00004ae9;
        11'h184: sin <= 32'h00004b19;
        11'h185: sin <= 32'h00004b49;
        11'h186: sin <= 32'h00004b79;
        11'h187: sin <= 32'h00004ba9;
        11'h188: sin <= 32'h00004bd9;
        11'h189: sin <= 32'h00004c09;
        11'h18a: sin <= 32'h00004c39;
        11'h18b: sin <= 32'h00004c69;
        11'h18c: sin <= 32'h00004c99;
        11'h18d: sin <= 32'h00004cc9;
        11'h18e: sin <= 32'h00004cf9;
        11'h18f: sin <= 32'h00004d29;
        11'h190: sin <= 32'h00004d59;
        11'h191: sin <= 32'h00004d89;
        11'h192: sin <= 32'h00004db9;
        11'h193: sin <= 32'h00004de8;
        11'h194: sin <= 32'h00004e18;
        11'h195: sin <= 32'h00004e48;
        11'h196: sin <= 32'h00004e78;
        11'h197: sin <= 32'h00004ea8;
        11'h198: sin <= 32'h00004ed8;
        11'h199: sin <= 32'h00004f08;
        11'h19a: sin <= 32'h00004f38;
        11'h19b: sin <= 32'h00004f67;
        11'h19c: sin <= 32'h00004f97;
        11'h19d: sin <= 32'h00004fc7;
        11'h19e: sin <= 32'h00004ff7;
        11'h19f: sin <= 32'h00005026;
        11'h1a0: sin <= 32'h00005056;
        11'h1a1: sin <= 32'h00005086;
        11'h1a2: sin <= 32'h000050b6;
        11'h1a3: sin <= 32'h000050e5;
        11'h1a4: sin <= 32'h00005115;
        11'h1a5: sin <= 32'h00005145;
        11'h1a6: sin <= 32'h00005174;
        11'h1a7: sin <= 32'h000051a4;
        11'h1a8: sin <= 32'h000051d4;
        11'h1a9: sin <= 32'h00005203;
        11'h1aa: sin <= 32'h00005233;
        11'h1ab: sin <= 32'h00005263;
        11'h1ac: sin <= 32'h00005292;
        11'h1ad: sin <= 32'h000052c2;
        11'h1ae: sin <= 32'h000052f1;
        11'h1af: sin <= 32'h00005321;
        11'h1b0: sin <= 32'h00005351;
        11'h1b1: sin <= 32'h00005380;
        11'h1b2: sin <= 32'h000053b0;
        11'h1b3: sin <= 32'h000053df;
        11'h1b4: sin <= 32'h0000540f;
        11'h1b5: sin <= 32'h0000543e;
        11'h1b6: sin <= 32'h0000546e;
        11'h1b7: sin <= 32'h0000549d;
        11'h1b8: sin <= 32'h000054cd;
        11'h1b9: sin <= 32'h000054fc;
        11'h1ba: sin <= 32'h0000552b;
        11'h1bb: sin <= 32'h0000555b;
        11'h1bc: sin <= 32'h0000558a;
        11'h1bd: sin <= 32'h000055ba;
        11'h1be: sin <= 32'h000055e9;
        11'h1bf: sin <= 32'h00005618;
        11'h1c0: sin <= 32'h00005648;
        11'h1c1: sin <= 32'h00005677;
        11'h1c2: sin <= 32'h000056a6;
        11'h1c3: sin <= 32'h000056d6;
        11'h1c4: sin <= 32'h00005705;
        11'h1c5: sin <= 32'h00005734;
        11'h1c6: sin <= 32'h00005764;
        11'h1c7: sin <= 32'h00005793;
        11'h1c8: sin <= 32'h000057c2;
        11'h1c9: sin <= 32'h000057f1;
        11'h1ca: sin <= 32'h00005821;
        11'h1cb: sin <= 32'h00005850;
        11'h1cc: sin <= 32'h0000587f;
        11'h1cd: sin <= 32'h000058ae;
        11'h1ce: sin <= 32'h000058dd;
        11'h1cf: sin <= 32'h0000590d;
        11'h1d0: sin <= 32'h0000593c;
        11'h1d1: sin <= 32'h0000596b;
        11'h1d2: sin <= 32'h0000599a;
        11'h1d3: sin <= 32'h000059c9;
        11'h1d4: sin <= 32'h000059f8;
        11'h1d5: sin <= 32'h00005a27;
        11'h1d6: sin <= 32'h00005a56;
        11'h1d7: sin <= 32'h00005a85;
        11'h1d8: sin <= 32'h00005ab4;
        11'h1d9: sin <= 32'h00005ae3;
        11'h1da: sin <= 32'h00005b12;
        11'h1db: sin <= 32'h00005b41;
        11'h1dc: sin <= 32'h00005b70;
        11'h1dd: sin <= 32'h00005b9f;
        11'h1de: sin <= 32'h00005bce;
        11'h1df: sin <= 32'h00005bfd;
        11'h1e0: sin <= 32'h00005c2c;
        11'h1e1: sin <= 32'h00005c5b;
        11'h1e2: sin <= 32'h00005c8a;
        11'h1e3: sin <= 32'h00005cb9;
        11'h1e4: sin <= 32'h00005ce8;
        11'h1e5: sin <= 32'h00005d16;
        11'h1e6: sin <= 32'h00005d45;
        11'h1e7: sin <= 32'h00005d74;
        11'h1e8: sin <= 32'h00005da3;
        11'h1e9: sin <= 32'h00005dd2;
        11'h1ea: sin <= 32'h00005e01;
        11'h1eb: sin <= 32'h00005e2f;
        11'h1ec: sin <= 32'h00005e5e;
        11'h1ed: sin <= 32'h00005e8d;
        11'h1ee: sin <= 32'h00005ebc;
        11'h1ef: sin <= 32'h00005eea;
        11'h1f0: sin <= 32'h00005f19;
        11'h1f1: sin <= 32'h00005f48;
        11'h1f2: sin <= 32'h00005f76;
        11'h1f3: sin <= 32'h00005fa5;
        11'h1f4: sin <= 32'h00005fd4;
        11'h1f5: sin <= 32'h00006002;
        11'h1f6: sin <= 32'h00006031;
        11'h1f7: sin <= 32'h0000605f;
        11'h1f8: sin <= 32'h0000608e;
        11'h1f9: sin <= 32'h000060bd;
        11'h1fa: sin <= 32'h000060eb;
        11'h1fb: sin <= 32'h0000611a;
        11'h1fc: sin <= 32'h00006148;
        11'h1fd: sin <= 32'h00006177;
        11'h1fe: sin <= 32'h000061a5;
        11'h1ff: sin <= 32'h000061d4;
        11'h200: sin <= 32'h00006202;
        11'h201: sin <= 32'h00006231;
        11'h202: sin <= 32'h0000625f;
        11'h203: sin <= 32'h0000628d;
        11'h204: sin <= 32'h000062bc;
        11'h205: sin <= 32'h000062ea;
        11'h206: sin <= 32'h00006319;
        11'h207: sin <= 32'h00006347;
        11'h208: sin <= 32'h00006375;
        11'h209: sin <= 32'h000063a4;
        11'h20a: sin <= 32'h000063d2;
        11'h20b: sin <= 32'h00006400;
        11'h20c: sin <= 32'h0000642e;
        11'h20d: sin <= 32'h0000645d;
        11'h20e: sin <= 32'h0000648b;
        11'h20f: sin <= 32'h000064b9;
        11'h210: sin <= 32'h000064e7;
        11'h211: sin <= 32'h00006516;
        11'h212: sin <= 32'h00006544;
        11'h213: sin <= 32'h00006572;
        11'h214: sin <= 32'h000065a0;
        11'h215: sin <= 32'h000065ce;
        11'h216: sin <= 32'h000065fd;
        11'h217: sin <= 32'h0000662b;
        11'h218: sin <= 32'h00006659;
        11'h219: sin <= 32'h00006687;
        11'h21a: sin <= 32'h000066b5;
        11'h21b: sin <= 32'h000066e3;
        11'h21c: sin <= 32'h00006711;
        11'h21d: sin <= 32'h0000673f;
        11'h21e: sin <= 32'h0000676d;
        11'h21f: sin <= 32'h0000679b;
        11'h220: sin <= 32'h000067c9;
        11'h221: sin <= 32'h000067f7;
        11'h222: sin <= 32'h00006825;
        11'h223: sin <= 32'h00006853;
        11'h224: sin <= 32'h00006881;
        11'h225: sin <= 32'h000068af;
        11'h226: sin <= 32'h000068dd;
        11'h227: sin <= 32'h0000690a;
        11'h228: sin <= 32'h00006938;
        11'h229: sin <= 32'h00006966;
        11'h22a: sin <= 32'h00006994;
        11'h22b: sin <= 32'h000069c2;
        11'h22c: sin <= 32'h000069ef;
        11'h22d: sin <= 32'h00006a1d;
        11'h22e: sin <= 32'h00006a4b;
        11'h22f: sin <= 32'h00006a79;
        11'h230: sin <= 32'h00006aa6;
        11'h231: sin <= 32'h00006ad4;
        11'h232: sin <= 32'h00006b02;
        11'h233: sin <= 32'h00006b30;
        11'h234: sin <= 32'h00006b5d;
        11'h235: sin <= 32'h00006b8b;
        11'h236: sin <= 32'h00006bb8;
        11'h237: sin <= 32'h00006be6;
        11'h238: sin <= 32'h00006c14;
        11'h239: sin <= 32'h00006c41;
        11'h23a: sin <= 32'h00006c6f;
        11'h23b: sin <= 32'h00006c9c;
        11'h23c: sin <= 32'h00006cca;
        11'h23d: sin <= 32'h00006cf7;
        11'h23e: sin <= 32'h00006d25;
        11'h23f: sin <= 32'h00006d52;
        11'h240: sin <= 32'h00006d80;
        11'h241: sin <= 32'h00006dad;
        11'h242: sin <= 32'h00006ddb;
        11'h243: sin <= 32'h00006e08;
        11'h244: sin <= 32'h00006e36;
        11'h245: sin <= 32'h00006e63;
        11'h246: sin <= 32'h00006e90;
        11'h247: sin <= 32'h00006ebe;
        11'h248: sin <= 32'h00006eeb;
        11'h249: sin <= 32'h00006f18;
        11'h24a: sin <= 32'h00006f46;
        11'h24b: sin <= 32'h00006f73;
        11'h24c: sin <= 32'h00006fa0;
        11'h24d: sin <= 32'h00006fcd;
        11'h24e: sin <= 32'h00006ffb;
        11'h24f: sin <= 32'h00007028;
        11'h250: sin <= 32'h00007055;
        11'h251: sin <= 32'h00007082;
        11'h252: sin <= 32'h000070af;
        11'h253: sin <= 32'h000070dd;
        11'h254: sin <= 32'h0000710a;
        11'h255: sin <= 32'h00007137;
        11'h256: sin <= 32'h00007164;
        11'h257: sin <= 32'h00007191;
        11'h258: sin <= 32'h000071be;
        11'h259: sin <= 32'h000071eb;
        11'h25a: sin <= 32'h00007218;
        11'h25b: sin <= 32'h00007245;
        11'h25c: sin <= 32'h00007272;
        11'h25d: sin <= 32'h0000729f;
        11'h25e: sin <= 32'h000072cc;
        11'h25f: sin <= 32'h000072f9;
        11'h260: sin <= 32'h00007326;
        11'h261: sin <= 32'h00007353;
        11'h262: sin <= 32'h00007380;
        11'h263: sin <= 32'h000073ad;
        11'h264: sin <= 32'h000073d9;
        11'h265: sin <= 32'h00007406;
        11'h266: sin <= 32'h00007433;
        11'h267: sin <= 32'h00007460;
        11'h268: sin <= 32'h0000748d;
        11'h269: sin <= 32'h000074b9;
        11'h26a: sin <= 32'h000074e6;
        11'h26b: sin <= 32'h00007513;
        11'h26c: sin <= 32'h00007540;
        11'h26d: sin <= 32'h0000756c;
        11'h26e: sin <= 32'h00007599;
        11'h26f: sin <= 32'h000075c6;
        11'h270: sin <= 32'h000075f2;
        11'h271: sin <= 32'h0000761f;
        11'h272: sin <= 32'h0000764b;
        11'h273: sin <= 32'h00007678;
        11'h274: sin <= 32'h000076a5;
        11'h275: sin <= 32'h000076d1;
        11'h276: sin <= 32'h000076fe;
        11'h277: sin <= 32'h0000772a;
        11'h278: sin <= 32'h00007757;
        11'h279: sin <= 32'h00007783;
        11'h27a: sin <= 32'h000077b0;
        11'h27b: sin <= 32'h000077dc;
        11'h27c: sin <= 32'h00007809;
        11'h27d: sin <= 32'h00007835;
        11'h27e: sin <= 32'h00007861;
        11'h27f: sin <= 32'h0000788e;
        11'h280: sin <= 32'h000078ba;
        11'h281: sin <= 32'h000078e6;
        11'h282: sin <= 32'h00007913;
        11'h283: sin <= 32'h0000793f;
        11'h284: sin <= 32'h0000796b;
        11'h285: sin <= 32'h00007998;
        11'h286: sin <= 32'h000079c4;
        11'h287: sin <= 32'h000079f0;
        11'h288: sin <= 32'h00007a1c;
        11'h289: sin <= 32'h00007a48;
        11'h28a: sin <= 32'h00007a75;
        11'h28b: sin <= 32'h00007aa1;
        11'h28c: sin <= 32'h00007acd;
        11'h28d: sin <= 32'h00007af9;
        11'h28e: sin <= 32'h00007b25;
        11'h28f: sin <= 32'h00007b51;
        11'h290: sin <= 32'h00007b7d;
        11'h291: sin <= 32'h00007ba9;
        11'h292: sin <= 32'h00007bd5;
        11'h293: sin <= 32'h00007c01;
        11'h294: sin <= 32'h00007c2d;
        11'h295: sin <= 32'h00007c59;
        11'h296: sin <= 32'h00007c85;
        11'h297: sin <= 32'h00007cb1;
        11'h298: sin <= 32'h00007cdd;
        11'h299: sin <= 32'h00007d09;
        11'h29a: sin <= 32'h00007d35;
        11'h29b: sin <= 32'h00007d61;
        11'h29c: sin <= 32'h00007d8c;
        11'h29d: sin <= 32'h00007db8;
        11'h29e: sin <= 32'h00007de4;
        11'h29f: sin <= 32'h00007e10;
        11'h2a0: sin <= 32'h00007e3c;
        11'h2a1: sin <= 32'h00007e67;
        11'h2a2: sin <= 32'h00007e93;
        11'h2a3: sin <= 32'h00007ebf;
        11'h2a4: sin <= 32'h00007eea;
        11'h2a5: sin <= 32'h00007f16;
        11'h2a6: sin <= 32'h00007f42;
        11'h2a7: sin <= 32'h00007f6d;
        11'h2a8: sin <= 32'h00007f99;
        11'h2a9: sin <= 32'h00007fc5;
        11'h2aa: sin <= 32'h00007ff0;
        11'h2ab: sin <= 32'h0000801c;
        11'h2ac: sin <= 32'h00008047;
        11'h2ad: sin <= 32'h00008073;
        11'h2ae: sin <= 32'h0000809e;
        11'h2af: sin <= 32'h000080ca;
        11'h2b0: sin <= 32'h000080f5;
        11'h2b1: sin <= 32'h00008121;
        11'h2b2: sin <= 32'h0000814c;
        11'h2b3: sin <= 32'h00008177;
        11'h2b4: sin <= 32'h000081a3;
        11'h2b5: sin <= 32'h000081ce;
        11'h2b6: sin <= 32'h000081f9;
        11'h2b7: sin <= 32'h00008225;
        11'h2b8: sin <= 32'h00008250;
        11'h2b9: sin <= 32'h0000827b;
        11'h2ba: sin <= 32'h000082a7;
        11'h2bb: sin <= 32'h000082d2;
        11'h2bc: sin <= 32'h000082fd;
        11'h2bd: sin <= 32'h00008328;
        11'h2be: sin <= 32'h00008353;
        11'h2bf: sin <= 32'h0000837f;
        11'h2c0: sin <= 32'h000083aa;
        11'h2c1: sin <= 32'h000083d5;
        11'h2c2: sin <= 32'h00008400;
        11'h2c3: sin <= 32'h0000842b;
        11'h2c4: sin <= 32'h00008456;
        11'h2c5: sin <= 32'h00008481;
        11'h2c6: sin <= 32'h000084ac;
        11'h2c7: sin <= 32'h000084d7;
        11'h2c8: sin <= 32'h00008502;
        11'h2c9: sin <= 32'h0000852d;
        11'h2ca: sin <= 32'h00008558;
        11'h2cb: sin <= 32'h00008583;
        11'h2cc: sin <= 32'h000085ae;
        11'h2cd: sin <= 32'h000085d9;
        11'h2ce: sin <= 32'h00008604;
        11'h2cf: sin <= 32'h0000862e;
        11'h2d0: sin <= 32'h00008659;
        11'h2d1: sin <= 32'h00008684;
        11'h2d2: sin <= 32'h000086af;
        11'h2d3: sin <= 32'h000086da;
        11'h2d4: sin <= 32'h00008704;
        11'h2d5: sin <= 32'h0000872f;
        11'h2d6: sin <= 32'h0000875a;
        11'h2d7: sin <= 32'h00008784;
        11'h2d8: sin <= 32'h000087af;
        11'h2d9: sin <= 32'h000087da;
        11'h2da: sin <= 32'h00008804;
        11'h2db: sin <= 32'h0000882f;
        11'h2dc: sin <= 32'h00008859;
        11'h2dd: sin <= 32'h00008884;
        11'h2de: sin <= 32'h000088ae;
        11'h2df: sin <= 32'h000088d9;
        11'h2e0: sin <= 32'h00008903;
        11'h2e1: sin <= 32'h0000892e;
        11'h2e2: sin <= 32'h00008958;
        11'h2e3: sin <= 32'h00008983;
        11'h2e4: sin <= 32'h000089ad;
        11'h2e5: sin <= 32'h000089d8;
        11'h2e6: sin <= 32'h00008a02;
        11'h2e7: sin <= 32'h00008a2c;
        11'h2e8: sin <= 32'h00008a57;
        11'h2e9: sin <= 32'h00008a81;
        11'h2ea: sin <= 32'h00008aab;
        11'h2eb: sin <= 32'h00008ad5;
        11'h2ec: sin <= 32'h00008b00;
        11'h2ed: sin <= 32'h00008b2a;
        11'h2ee: sin <= 32'h00008b54;
        11'h2ef: sin <= 32'h00008b7e;
        11'h2f0: sin <= 32'h00008ba8;
        11'h2f1: sin <= 32'h00008bd3;
        11'h2f2: sin <= 32'h00008bfd;
        11'h2f3: sin <= 32'h00008c27;
        11'h2f4: sin <= 32'h00008c51;
        11'h2f5: sin <= 32'h00008c7b;
        11'h2f6: sin <= 32'h00008ca5;
        11'h2f7: sin <= 32'h00008ccf;
        11'h2f8: sin <= 32'h00008cf9;
        11'h2f9: sin <= 32'h00008d23;
        11'h2fa: sin <= 32'h00008d4d;
        11'h2fb: sin <= 32'h00008d77;
        11'h2fc: sin <= 32'h00008da1;
        11'h2fd: sin <= 32'h00008dcb;
        11'h2fe: sin <= 32'h00008df4;
        11'h2ff: sin <= 32'h00008e1e;
        11'h300: sin <= 32'h00008e48;
        11'h301: sin <= 32'h00008e72;
        11'h302: sin <= 32'h00008e9c;
        11'h303: sin <= 32'h00008ec5;
        11'h304: sin <= 32'h00008eef;
        11'h305: sin <= 32'h00008f19;
        11'h306: sin <= 32'h00008f43;
        11'h307: sin <= 32'h00008f6c;
        11'h308: sin <= 32'h00008f96;
        11'h309: sin <= 32'h00008fbf;
        11'h30a: sin <= 32'h00008fe9;
        11'h30b: sin <= 32'h00009013;
        11'h30c: sin <= 32'h0000903c;
        11'h30d: sin <= 32'h00009066;
        11'h30e: sin <= 32'h0000908f;
        11'h30f: sin <= 32'h000090b9;
        11'h310: sin <= 32'h000090e2;
        11'h311: sin <= 32'h0000910c;
        11'h312: sin <= 32'h00009135;
        11'h313: sin <= 32'h0000915f;
        11'h314: sin <= 32'h00009188;
        11'h315: sin <= 32'h000091b1;
        11'h316: sin <= 32'h000091db;
        11'h317: sin <= 32'h00009204;
        11'h318: sin <= 32'h0000922d;
        11'h319: sin <= 32'h00009256;
        11'h31a: sin <= 32'h00009280;
        11'h31b: sin <= 32'h000092a9;
        11'h31c: sin <= 32'h000092d2;
        11'h31d: sin <= 32'h000092fb;
        11'h31e: sin <= 32'h00009324;
        11'h31f: sin <= 32'h0000934e;
        11'h320: sin <= 32'h00009377;
        11'h321: sin <= 32'h000093a0;
        11'h322: sin <= 32'h000093c9;
        11'h323: sin <= 32'h000093f2;
        11'h324: sin <= 32'h0000941b;
        11'h325: sin <= 32'h00009444;
        11'h326: sin <= 32'h0000946d;
        11'h327: sin <= 32'h00009496;
        11'h328: sin <= 32'h000094bf;
        11'h329: sin <= 32'h000094e8;
        11'h32a: sin <= 32'h00009511;
        11'h32b: sin <= 32'h0000953a;
        11'h32c: sin <= 32'h00009562;
        11'h32d: sin <= 32'h0000958b;
        11'h32e: sin <= 32'h000095b4;
        11'h32f: sin <= 32'h000095dd;
        11'h330: sin <= 32'h00009606;
        11'h331: sin <= 32'h0000962e;
        11'h332: sin <= 32'h00009657;
        11'h333: sin <= 32'h00009680;
        11'h334: sin <= 32'h000096a8;
        11'h335: sin <= 32'h000096d1;
        11'h336: sin <= 32'h000096fa;
        11'h337: sin <= 32'h00009722;
        11'h338: sin <= 32'h0000974b;
        11'h339: sin <= 32'h00009773;
        11'h33a: sin <= 32'h0000979c;
        11'h33b: sin <= 32'h000097c4;
        11'h33c: sin <= 32'h000097ed;
        11'h33d: sin <= 32'h00009815;
        11'h33e: sin <= 32'h0000983e;
        11'h33f: sin <= 32'h00009866;
        11'h340: sin <= 32'h0000988f;
        11'h341: sin <= 32'h000098b7;
        11'h342: sin <= 32'h000098df;
        11'h343: sin <= 32'h00009908;
        11'h344: sin <= 32'h00009930;
        11'h345: sin <= 32'h00009958;
        11'h346: sin <= 32'h00009981;
        11'h347: sin <= 32'h000099a9;
        11'h348: sin <= 32'h000099d1;
        11'h349: sin <= 32'h000099f9;
        11'h34a: sin <= 32'h00009a21;
        11'h34b: sin <= 32'h00009a49;
        11'h34c: sin <= 32'h00009a72;
        11'h34d: sin <= 32'h00009a9a;
        11'h34e: sin <= 32'h00009ac2;
        11'h34f: sin <= 32'h00009aea;
        11'h350: sin <= 32'h00009b12;
        11'h351: sin <= 32'h00009b3a;
        11'h352: sin <= 32'h00009b62;
        11'h353: sin <= 32'h00009b8a;
        11'h354: sin <= 32'h00009bb2;
        11'h355: sin <= 32'h00009bda;
        11'h356: sin <= 32'h00009c01;
        11'h357: sin <= 32'h00009c29;
        11'h358: sin <= 32'h00009c51;
        11'h359: sin <= 32'h00009c79;
        11'h35a: sin <= 32'h00009ca1;
        11'h35b: sin <= 32'h00009cc9;
        11'h35c: sin <= 32'h00009cf0;
        11'h35d: sin <= 32'h00009d18;
        11'h35e: sin <= 32'h00009d40;
        11'h35f: sin <= 32'h00009d67;
        11'h360: sin <= 32'h00009d8f;
        11'h361: sin <= 32'h00009db7;
        11'h362: sin <= 32'h00009dde;
        11'h363: sin <= 32'h00009e06;
        11'h364: sin <= 32'h00009e2d;
        11'h365: sin <= 32'h00009e55;
        11'h366: sin <= 32'h00009e7c;
        11'h367: sin <= 32'h00009ea4;
        11'h368: sin <= 32'h00009ecb;
        11'h369: sin <= 32'h00009ef3;
        11'h36a: sin <= 32'h00009f1a;
        11'h36b: sin <= 32'h00009f42;
        11'h36c: sin <= 32'h00009f69;
        11'h36d: sin <= 32'h00009f90;
        11'h36e: sin <= 32'h00009fb8;
        11'h36f: sin <= 32'h00009fdf;
        11'h370: sin <= 32'h0000a006;
        11'h371: sin <= 32'h0000a02d;
        11'h372: sin <= 32'h0000a055;
        11'h373: sin <= 32'h0000a07c;
        11'h374: sin <= 32'h0000a0a3;
        11'h375: sin <= 32'h0000a0ca;
        11'h376: sin <= 32'h0000a0f1;
        11'h377: sin <= 32'h0000a118;
        11'h378: sin <= 32'h0000a13f;
        11'h379: sin <= 32'h0000a166;
        11'h37a: sin <= 32'h0000a18d;
        11'h37b: sin <= 32'h0000a1b4;
        11'h37c: sin <= 32'h0000a1db;
        11'h37d: sin <= 32'h0000a202;
        11'h37e: sin <= 32'h0000a229;
        11'h37f: sin <= 32'h0000a250;
        11'h380: sin <= 32'h0000a277;
        11'h381: sin <= 32'h0000a29e;
        11'h382: sin <= 32'h0000a2c5;
        11'h383: sin <= 32'h0000a2ec;
        11'h384: sin <= 32'h0000a312;
        11'h385: sin <= 32'h0000a339;
        11'h386: sin <= 32'h0000a360;
        11'h387: sin <= 32'h0000a386;
        11'h388: sin <= 32'h0000a3ad;
        11'h389: sin <= 32'h0000a3d4;
        11'h38a: sin <= 32'h0000a3fa;
        11'h38b: sin <= 32'h0000a421;
        11'h38c: sin <= 32'h0000a448;
        11'h38d: sin <= 32'h0000a46e;
        11'h38e: sin <= 32'h0000a495;
        11'h38f: sin <= 32'h0000a4bb;
        11'h390: sin <= 32'h0000a4e2;
        11'h391: sin <= 32'h0000a508;
        11'h392: sin <= 32'h0000a52f;
        11'h393: sin <= 32'h0000a555;
        11'h394: sin <= 32'h0000a57b;
        11'h395: sin <= 32'h0000a5a2;
        11'h396: sin <= 32'h0000a5c8;
        11'h397: sin <= 32'h0000a5ee;
        11'h398: sin <= 32'h0000a615;
        11'h399: sin <= 32'h0000a63b;
        11'h39a: sin <= 32'h0000a661;
        11'h39b: sin <= 32'h0000a687;
        11'h39c: sin <= 32'h0000a6ae;
        11'h39d: sin <= 32'h0000a6d4;
        11'h39e: sin <= 32'h0000a6fa;
        11'h39f: sin <= 32'h0000a720;
        11'h3a0: sin <= 32'h0000a746;
        11'h3a1: sin <= 32'h0000a76c;
        11'h3a2: sin <= 32'h0000a792;
        11'h3a3: sin <= 32'h0000a7b8;
        11'h3a4: sin <= 32'h0000a7de;
        11'h3a5: sin <= 32'h0000a804;
        11'h3a6: sin <= 32'h0000a82a;
        11'h3a7: sin <= 32'h0000a850;
        11'h3a8: sin <= 32'h0000a876;
        11'h3a9: sin <= 32'h0000a89c;
        11'h3aa: sin <= 32'h0000a8c1;
        11'h3ab: sin <= 32'h0000a8e7;
        11'h3ac: sin <= 32'h0000a90d;
        11'h3ad: sin <= 32'h0000a933;
        11'h3ae: sin <= 32'h0000a958;
        11'h3af: sin <= 32'h0000a97e;
        11'h3b0: sin <= 32'h0000a9a4;
        11'h3b1: sin <= 32'h0000a9c9;
        11'h3b2: sin <= 32'h0000a9ef;
        11'h3b3: sin <= 32'h0000aa15;
        11'h3b4: sin <= 32'h0000aa3a;
        11'h3b5: sin <= 32'h0000aa60;
        11'h3b6: sin <= 32'h0000aa85;
        11'h3b7: sin <= 32'h0000aaab;
        11'h3b8: sin <= 32'h0000aad0;
        11'h3b9: sin <= 32'h0000aaf6;
        11'h3ba: sin <= 32'h0000ab1b;
        11'h3bb: sin <= 32'h0000ab41;
        11'h3bc: sin <= 32'h0000ab66;
        11'h3bd: sin <= 32'h0000ab8b;
        11'h3be: sin <= 32'h0000abb1;
        11'h3bf: sin <= 32'h0000abd6;
        11'h3c0: sin <= 32'h0000abfb;
        11'h3c1: sin <= 32'h0000ac20;
        11'h3c2: sin <= 32'h0000ac46;
        11'h3c3: sin <= 32'h0000ac6b;
        11'h3c4: sin <= 32'h0000ac90;
        11'h3c5: sin <= 32'h0000acb5;
        11'h3c6: sin <= 32'h0000acda;
        11'h3c7: sin <= 32'h0000acff;
        11'h3c8: sin <= 32'h0000ad24;
        11'h3c9: sin <= 32'h0000ad49;
        11'h3ca: sin <= 32'h0000ad6e;
        11'h3cb: sin <= 32'h0000ad93;
        11'h3cc: sin <= 32'h0000adb8;
        11'h3cd: sin <= 32'h0000addd;
        11'h3ce: sin <= 32'h0000ae02;
        11'h3cf: sin <= 32'h0000ae27;
        11'h3d0: sin <= 32'h0000ae4c;
        11'h3d1: sin <= 32'h0000ae71;
        11'h3d2: sin <= 32'h0000ae95;
        11'h3d3: sin <= 32'h0000aeba;
        11'h3d4: sin <= 32'h0000aedf;
        11'h3d5: sin <= 32'h0000af04;
        11'h3d6: sin <= 32'h0000af28;
        11'h3d7: sin <= 32'h0000af4d;
        11'h3d8: sin <= 32'h0000af72;
        11'h3d9: sin <= 32'h0000af96;
        11'h3da: sin <= 32'h0000afbb;
        11'h3db: sin <= 32'h0000afdf;
        11'h3dc: sin <= 32'h0000b004;
        11'h3dd: sin <= 32'h0000b028;
        11'h3de: sin <= 32'h0000b04d;
        11'h3df: sin <= 32'h0000b071;
        11'h3e0: sin <= 32'h0000b096;
        11'h3e1: sin <= 32'h0000b0ba;
        11'h3e2: sin <= 32'h0000b0de;
        11'h3e3: sin <= 32'h0000b103;
        11'h3e4: sin <= 32'h0000b127;
        11'h3e5: sin <= 32'h0000b14b;
        11'h3e6: sin <= 32'h0000b170;
        11'h3e7: sin <= 32'h0000b194;
        11'h3e8: sin <= 32'h0000b1b8;
        11'h3e9: sin <= 32'h0000b1dc;
        11'h3ea: sin <= 32'h0000b200;
        11'h3eb: sin <= 32'h0000b225;
        11'h3ec: sin <= 32'h0000b249;
        11'h3ed: sin <= 32'h0000b26d;
        11'h3ee: sin <= 32'h0000b291;
        11'h3ef: sin <= 32'h0000b2b5;
        11'h3f0: sin <= 32'h0000b2d9;
        11'h3f1: sin <= 32'h0000b2fd;
        11'h3f2: sin <= 32'h0000b321;
        11'h3f3: sin <= 32'h0000b345;
        11'h3f4: sin <= 32'h0000b369;
        11'h3f5: sin <= 32'h0000b38c;
        11'h3f6: sin <= 32'h0000b3b0;
        11'h3f7: sin <= 32'h0000b3d4;
        11'h3f8: sin <= 32'h0000b3f8;
        11'h3f9: sin <= 32'h0000b41c;
        11'h3fa: sin <= 32'h0000b43f;
        11'h3fb: sin <= 32'h0000b463;
        11'h3fc: sin <= 32'h0000b487;
        11'h3fd: sin <= 32'h0000b4aa;
        11'h3fe: sin <= 32'h0000b4ce;
        11'h3ff: sin <= 32'h0000b4f1;
        11'h400: sin <= 32'h0000b515;
        11'h401: sin <= 32'h0000b539;
        11'h402: sin <= 32'h0000b55c;
        11'h403: sin <= 32'h0000b580;
        11'h404: sin <= 32'h0000b5a3;
        11'h405: sin <= 32'h0000b5c6;
        11'h406: sin <= 32'h0000b5ea;
        11'h407: sin <= 32'h0000b60d;
        11'h408: sin <= 32'h0000b631;
        11'h409: sin <= 32'h0000b654;
        11'h40a: sin <= 32'h0000b677;
        11'h40b: sin <= 32'h0000b69a;
        11'h40c: sin <= 32'h0000b6be;
        11'h40d: sin <= 32'h0000b6e1;
        11'h40e: sin <= 32'h0000b704;
        11'h40f: sin <= 32'h0000b727;
        11'h410: sin <= 32'h0000b74a;
        11'h411: sin <= 32'h0000b76d;
        11'h412: sin <= 32'h0000b790;
        11'h413: sin <= 32'h0000b7b3;
        11'h414: sin <= 32'h0000b7d6;
        11'h415: sin <= 32'h0000b7f9;
        11'h416: sin <= 32'h0000b81c;
        11'h417: sin <= 32'h0000b83f;
        11'h418: sin <= 32'h0000b862;
        11'h419: sin <= 32'h0000b885;
        11'h41a: sin <= 32'h0000b8a8;
        11'h41b: sin <= 32'h0000b8cb;
        11'h41c: sin <= 32'h0000b8ee;
        11'h41d: sin <= 32'h0000b910;
        11'h41e: sin <= 32'h0000b933;
        11'h41f: sin <= 32'h0000b956;
        11'h420: sin <= 32'h0000b978;
        11'h421: sin <= 32'h0000b99b;
        11'h422: sin <= 32'h0000b9be;
        11'h423: sin <= 32'h0000b9e0;
        11'h424: sin <= 32'h0000ba03;
        11'h425: sin <= 32'h0000ba25;
        11'h426: sin <= 32'h0000ba48;
        11'h427: sin <= 32'h0000ba6a;
        11'h428: sin <= 32'h0000ba8d;
        11'h429: sin <= 32'h0000baaf;
        11'h42a: sin <= 32'h0000bad2;
        11'h42b: sin <= 32'h0000baf4;
        11'h42c: sin <= 32'h0000bb16;
        11'h42d: sin <= 32'h0000bb39;
        11'h42e: sin <= 32'h0000bb5b;
        11'h42f: sin <= 32'h0000bb7d;
        11'h430: sin <= 32'h0000bb9f;
        11'h431: sin <= 32'h0000bbc2;
        11'h432: sin <= 32'h0000bbe4;
        11'h433: sin <= 32'h0000bc06;
        11'h434: sin <= 32'h0000bc28;
        11'h435: sin <= 32'h0000bc4a;
        11'h436: sin <= 32'h0000bc6c;
        11'h437: sin <= 32'h0000bc8e;
        11'h438: sin <= 32'h0000bcb0;
        11'h439: sin <= 32'h0000bcd2;
        11'h43a: sin <= 32'h0000bcf4;
        11'h43b: sin <= 32'h0000bd16;
        11'h43c: sin <= 32'h0000bd38;
        11'h43d: sin <= 32'h0000bd5a;
        11'h43e: sin <= 32'h0000bd7c;
        11'h43f: sin <= 32'h0000bd9d;
        11'h440: sin <= 32'h0000bdbf;
        11'h441: sin <= 32'h0000bde1;
        11'h442: sin <= 32'h0000be03;
        11'h443: sin <= 32'h0000be24;
        11'h444: sin <= 32'h0000be46;
        11'h445: sin <= 32'h0000be68;
        11'h446: sin <= 32'h0000be89;
        11'h447: sin <= 32'h0000beab;
        11'h448: sin <= 32'h0000becc;
        11'h449: sin <= 32'h0000beee;
        11'h44a: sin <= 32'h0000bf0f;
        11'h44b: sin <= 32'h0000bf31;
        11'h44c: sin <= 32'h0000bf52;
        11'h44d: sin <= 32'h0000bf74;
        11'h44e: sin <= 32'h0000bf95;
        11'h44f: sin <= 32'h0000bfb6;
        11'h450: sin <= 32'h0000bfd8;
        11'h451: sin <= 32'h0000bff9;
        11'h452: sin <= 32'h0000c01a;
        11'h453: sin <= 32'h0000c03b;
        11'h454: sin <= 32'h0000c05d;
        11'h455: sin <= 32'h0000c07e;
        11'h456: sin <= 32'h0000c09f;
        11'h457: sin <= 32'h0000c0c0;
        11'h458: sin <= 32'h0000c0e1;
        11'h459: sin <= 32'h0000c102;
        11'h45a: sin <= 32'h0000c123;
        11'h45b: sin <= 32'h0000c144;
        11'h45c: sin <= 32'h0000c165;
        11'h45d: sin <= 32'h0000c186;
        11'h45e: sin <= 32'h0000c1a7;
        11'h45f: sin <= 32'h0000c1c8;
        11'h460: sin <= 32'h0000c1e9;
        11'h461: sin <= 32'h0000c209;
        11'h462: sin <= 32'h0000c22a;
        11'h463: sin <= 32'h0000c24b;
        11'h464: sin <= 32'h0000c26c;
        11'h465: sin <= 32'h0000c28c;
        11'h466: sin <= 32'h0000c2ad;
        11'h467: sin <= 32'h0000c2ce;
        11'h468: sin <= 32'h0000c2ee;
        11'h469: sin <= 32'h0000c30f;
        11'h46a: sin <= 32'h0000c32f;
        11'h46b: sin <= 32'h0000c350;
        11'h46c: sin <= 32'h0000c370;
        11'h46d: sin <= 32'h0000c391;
        11'h46e: sin <= 32'h0000c3b1;
        11'h46f: sin <= 32'h0000c3d2;
        11'h470: sin <= 32'h0000c3f2;
        11'h471: sin <= 32'h0000c413;
        11'h472: sin <= 32'h0000c433;
        11'h473: sin <= 32'h0000c453;
        11'h474: sin <= 32'h0000c473;
        11'h475: sin <= 32'h0000c494;
        11'h476: sin <= 32'h0000c4b4;
        11'h477: sin <= 32'h0000c4d4;
        11'h478: sin <= 32'h0000c4f4;
        11'h479: sin <= 32'h0000c514;
        11'h47a: sin <= 32'h0000c534;
        11'h47b: sin <= 32'h0000c554;
        11'h47c: sin <= 32'h0000c574;
        11'h47d: sin <= 32'h0000c594;
        11'h47e: sin <= 32'h0000c5b4;
        11'h47f: sin <= 32'h0000c5d4;
        11'h480: sin <= 32'h0000c5f4;
        11'h481: sin <= 32'h0000c614;
        11'h482: sin <= 32'h0000c634;
        11'h483: sin <= 32'h0000c654;
        11'h484: sin <= 32'h0000c673;
        11'h485: sin <= 32'h0000c693;
        11'h486: sin <= 32'h0000c6b3;
        11'h487: sin <= 32'h0000c6d3;
        11'h488: sin <= 32'h0000c6f2;
        11'h489: sin <= 32'h0000c712;
        11'h48a: sin <= 32'h0000c732;
        11'h48b: sin <= 32'h0000c751;
        11'h48c: sin <= 32'h0000c771;
        11'h48d: sin <= 32'h0000c790;
        11'h48e: sin <= 32'h0000c7b0;
        11'h48f: sin <= 32'h0000c7cf;
        11'h490: sin <= 32'h0000c7ef;
        11'h491: sin <= 32'h0000c80e;
        11'h492: sin <= 32'h0000c82d;
        11'h493: sin <= 32'h0000c84d;
        11'h494: sin <= 32'h0000c86c;
        11'h495: sin <= 32'h0000c88b;
        11'h496: sin <= 32'h0000c8aa;
        11'h497: sin <= 32'h0000c8ca;
        11'h498: sin <= 32'h0000c8e9;
        11'h499: sin <= 32'h0000c908;
        11'h49a: sin <= 32'h0000c927;
        11'h49b: sin <= 32'h0000c946;
        11'h49c: sin <= 32'h0000c965;
        11'h49d: sin <= 32'h0000c984;
        11'h49e: sin <= 32'h0000c9a3;
        11'h49f: sin <= 32'h0000c9c2;
        11'h4a0: sin <= 32'h0000c9e1;
        11'h4a1: sin <= 32'h0000ca00;
        11'h4a2: sin <= 32'h0000ca1f;
        11'h4a3: sin <= 32'h0000ca3e;
        11'h4a4: sin <= 32'h0000ca5d;
        11'h4a5: sin <= 32'h0000ca7b;
        11'h4a6: sin <= 32'h0000ca9a;
        11'h4a7: sin <= 32'h0000cab9;
        11'h4a8: sin <= 32'h0000cad8;
        11'h4a9: sin <= 32'h0000caf6;
        11'h4aa: sin <= 32'h0000cb15;
        11'h4ab: sin <= 32'h0000cb33;
        11'h4ac: sin <= 32'h0000cb52;
        11'h4ad: sin <= 32'h0000cb71;
        11'h4ae: sin <= 32'h0000cb8f;
        11'h4af: sin <= 32'h0000cbae;
        11'h4b0: sin <= 32'h0000cbcc;
        11'h4b1: sin <= 32'h0000cbea;
        11'h4b2: sin <= 32'h0000cc09;
        11'h4b3: sin <= 32'h0000cc27;
        11'h4b4: sin <= 32'h0000cc45;
        11'h4b5: sin <= 32'h0000cc64;
        11'h4b6: sin <= 32'h0000cc82;
        11'h4b7: sin <= 32'h0000cca0;
        11'h4b8: sin <= 32'h0000ccbe;
        11'h4b9: sin <= 32'h0000ccdd;
        11'h4ba: sin <= 32'h0000ccfb;
        11'h4bb: sin <= 32'h0000cd19;
        11'h4bc: sin <= 32'h0000cd37;
        11'h4bd: sin <= 32'h0000cd55;
        11'h4be: sin <= 32'h0000cd73;
        11'h4bf: sin <= 32'h0000cd91;
        11'h4c0: sin <= 32'h0000cdaf;
        11'h4c1: sin <= 32'h0000cdcd;
        11'h4c2: sin <= 32'h0000cdeb;
        11'h4c3: sin <= 32'h0000ce09;
        11'h4c4: sin <= 32'h0000ce26;
        11'h4c5: sin <= 32'h0000ce44;
        11'h4c6: sin <= 32'h0000ce62;
        11'h4c7: sin <= 32'h0000ce80;
        11'h4c8: sin <= 32'h0000ce9d;
        11'h4c9: sin <= 32'h0000cebb;
        11'h4ca: sin <= 32'h0000ced9;
        11'h4cb: sin <= 32'h0000cef6;
        11'h4cc: sin <= 32'h0000cf14;
        11'h4cd: sin <= 32'h0000cf32;
        11'h4ce: sin <= 32'h0000cf4f;
        11'h4cf: sin <= 32'h0000cf6d;
        11'h4d0: sin <= 32'h0000cf8a;
        11'h4d1: sin <= 32'h0000cfa7;
        11'h4d2: sin <= 32'h0000cfc5;
        11'h4d3: sin <= 32'h0000cfe2;
        11'h4d4: sin <= 32'h0000d000;
        11'h4d5: sin <= 32'h0000d01d;
        11'h4d6: sin <= 32'h0000d03a;
        11'h4d7: sin <= 32'h0000d057;
        11'h4d8: sin <= 32'h0000d075;
        11'h4d9: sin <= 32'h0000d092;
        11'h4da: sin <= 32'h0000d0af;
        11'h4db: sin <= 32'h0000d0cc;
        11'h4dc: sin <= 32'h0000d0e9;
        11'h4dd: sin <= 32'h0000d106;
        11'h4de: sin <= 32'h0000d123;
        11'h4df: sin <= 32'h0000d140;
        11'h4e0: sin <= 32'h0000d15d;
        11'h4e1: sin <= 32'h0000d17a;
        11'h4e2: sin <= 32'h0000d197;
        11'h4e3: sin <= 32'h0000d1b4;
        11'h4e4: sin <= 32'h0000d1d1;
        11'h4e5: sin <= 32'h0000d1ed;
        11'h4e6: sin <= 32'h0000d20a;
        11'h4e7: sin <= 32'h0000d227;
        11'h4e8: sin <= 32'h0000d244;
        11'h4e9: sin <= 32'h0000d260;
        11'h4ea: sin <= 32'h0000d27d;
        11'h4eb: sin <= 32'h0000d299;
        11'h4ec: sin <= 32'h0000d2b6;
        11'h4ed: sin <= 32'h0000d2d3;
        11'h4ee: sin <= 32'h0000d2ef;
        11'h4ef: sin <= 32'h0000d30c;
        11'h4f0: sin <= 32'h0000d328;
        11'h4f1: sin <= 32'h0000d344;
        11'h4f2: sin <= 32'h0000d361;
        11'h4f3: sin <= 32'h0000d37d;
        11'h4f4: sin <= 32'h0000d399;
        11'h4f5: sin <= 32'h0000d3b6;
        11'h4f6: sin <= 32'h0000d3d2;
        11'h4f7: sin <= 32'h0000d3ee;
        11'h4f8: sin <= 32'h0000d40a;
        11'h4f9: sin <= 32'h0000d427;
        11'h4fa: sin <= 32'h0000d443;
        11'h4fb: sin <= 32'h0000d45f;
        11'h4fc: sin <= 32'h0000d47b;
        11'h4fd: sin <= 32'h0000d497;
        11'h4fe: sin <= 32'h0000d4b3;
        11'h4ff: sin <= 32'h0000d4cf;
        11'h500: sin <= 32'h0000d4eb;
        11'h501: sin <= 32'h0000d507;
        11'h502: sin <= 32'h0000d523;
        11'h503: sin <= 32'h0000d53e;
        11'h504: sin <= 32'h0000d55a;
        11'h505: sin <= 32'h0000d576;
        11'h506: sin <= 32'h0000d592;
        11'h507: sin <= 32'h0000d5ad;
        11'h508: sin <= 32'h0000d5c9;
        11'h509: sin <= 32'h0000d5e5;
        11'h50a: sin <= 32'h0000d600;
        11'h50b: sin <= 32'h0000d61c;
        11'h50c: sin <= 32'h0000d638;
        11'h50d: sin <= 32'h0000d653;
        11'h50e: sin <= 32'h0000d66f;
        11'h50f: sin <= 32'h0000d68a;
        11'h510: sin <= 32'h0000d6a5;
        11'h511: sin <= 32'h0000d6c1;
        11'h512: sin <= 32'h0000d6dc;
        11'h513: sin <= 32'h0000d6f7;
        11'h514: sin <= 32'h0000d713;
        11'h515: sin <= 32'h0000d72e;
        11'h516: sin <= 32'h0000d749;
        11'h517: sin <= 32'h0000d764;
        11'h518: sin <= 32'h0000d780;
        11'h519: sin <= 32'h0000d79b;
        11'h51a: sin <= 32'h0000d7b6;
        11'h51b: sin <= 32'h0000d7d1;
        11'h51c: sin <= 32'h0000d7ec;
        11'h51d: sin <= 32'h0000d807;
        11'h51e: sin <= 32'h0000d822;
        11'h51f: sin <= 32'h0000d83d;
        11'h520: sin <= 32'h0000d858;
        11'h521: sin <= 32'h0000d873;
        11'h522: sin <= 32'h0000d88d;
        11'h523: sin <= 32'h0000d8a8;
        11'h524: sin <= 32'h0000d8c3;
        11'h525: sin <= 32'h0000d8de;
        11'h526: sin <= 32'h0000d8f8;
        11'h527: sin <= 32'h0000d913;
        11'h528: sin <= 32'h0000d92e;
        11'h529: sin <= 32'h0000d948;
        11'h52a: sin <= 32'h0000d963;
        11'h52b: sin <= 32'h0000d97d;
        11'h52c: sin <= 32'h0000d998;
        11'h52d: sin <= 32'h0000d9b2;
        11'h52e: sin <= 32'h0000d9cd;
        11'h52f: sin <= 32'h0000d9e7;
        11'h530: sin <= 32'h0000da02;
        11'h531: sin <= 32'h0000da1c;
        11'h532: sin <= 32'h0000da36;
        11'h533: sin <= 32'h0000da51;
        11'h534: sin <= 32'h0000da6b;
        11'h535: sin <= 32'h0000da85;
        11'h536: sin <= 32'h0000da9f;
        11'h537: sin <= 32'h0000dab9;
        11'h538: sin <= 32'h0000dad3;
        11'h539: sin <= 32'h0000daee;
        11'h53a: sin <= 32'h0000db08;
        11'h53b: sin <= 32'h0000db22;
        11'h53c: sin <= 32'h0000db3c;
        11'h53d: sin <= 32'h0000db56;
        11'h53e: sin <= 32'h0000db6f;
        11'h53f: sin <= 32'h0000db89;
        11'h540: sin <= 32'h0000dba3;
        11'h541: sin <= 32'h0000dbbd;
        11'h542: sin <= 32'h0000dbd7;
        11'h543: sin <= 32'h0000dbf1;
        11'h544: sin <= 32'h0000dc0a;
        11'h545: sin <= 32'h0000dc24;
        11'h546: sin <= 32'h0000dc3e;
        11'h547: sin <= 32'h0000dc57;
        11'h548: sin <= 32'h0000dc71;
        11'h549: sin <= 32'h0000dc8a;
        11'h54a: sin <= 32'h0000dca4;
        11'h54b: sin <= 32'h0000dcbd;
        11'h54c: sin <= 32'h0000dcd7;
        11'h54d: sin <= 32'h0000dcf0;
        11'h54e: sin <= 32'h0000dd0a;
        11'h54f: sin <= 32'h0000dd23;
        11'h550: sin <= 32'h0000dd3c;
        11'h551: sin <= 32'h0000dd56;
        11'h552: sin <= 32'h0000dd6f;
        11'h553: sin <= 32'h0000dd88;
        11'h554: sin <= 32'h0000dda1;
        11'h555: sin <= 32'h0000ddba;
        11'h556: sin <= 32'h0000ddd3;
        11'h557: sin <= 32'h0000dded;
        11'h558: sin <= 32'h0000de06;
        11'h559: sin <= 32'h0000de1f;
        11'h55a: sin <= 32'h0000de38;
        11'h55b: sin <= 32'h0000de51;
        11'h55c: sin <= 32'h0000de69;
        11'h55d: sin <= 32'h0000de82;
        11'h55e: sin <= 32'h0000de9b;
        11'h55f: sin <= 32'h0000deb4;
        11'h560: sin <= 32'h0000decd;
        11'h561: sin <= 32'h0000dee6;
        11'h562: sin <= 32'h0000defe;
        11'h563: sin <= 32'h0000df17;
        11'h564: sin <= 32'h0000df30;
        11'h565: sin <= 32'h0000df48;
        11'h566: sin <= 32'h0000df61;
        11'h567: sin <= 32'h0000df79;
        11'h568: sin <= 32'h0000df92;
        11'h569: sin <= 32'h0000dfaa;
        11'h56a: sin <= 32'h0000dfc3;
        11'h56b: sin <= 32'h0000dfdb;
        11'h56c: sin <= 32'h0000dff4;
        11'h56d: sin <= 32'h0000e00c;
        11'h56e: sin <= 32'h0000e024;
        11'h56f: sin <= 32'h0000e03c;
        11'h570: sin <= 32'h0000e055;
        11'h571: sin <= 32'h0000e06d;
        11'h572: sin <= 32'h0000e085;
        11'h573: sin <= 32'h0000e09d;
        11'h574: sin <= 32'h0000e0b5;
        11'h575: sin <= 32'h0000e0cd;
        11'h576: sin <= 32'h0000e0e5;
        11'h577: sin <= 32'h0000e0fd;
        11'h578: sin <= 32'h0000e115;
        11'h579: sin <= 32'h0000e12d;
        11'h57a: sin <= 32'h0000e145;
        11'h57b: sin <= 32'h0000e15d;
        11'h57c: sin <= 32'h0000e175;
        11'h57d: sin <= 32'h0000e18d;
        11'h57e: sin <= 32'h0000e1a5;
        11'h57f: sin <= 32'h0000e1bc;
        11'h580: sin <= 32'h0000e1d4;
        11'h581: sin <= 32'h0000e1ec;
        11'h582: sin <= 32'h0000e203;
        11'h583: sin <= 32'h0000e21b;
        11'h584: sin <= 32'h0000e232;
        11'h585: sin <= 32'h0000e24a;
        11'h586: sin <= 32'h0000e261;
        11'h587: sin <= 32'h0000e279;
        11'h588: sin <= 32'h0000e290;
        11'h589: sin <= 32'h0000e2a8;
        11'h58a: sin <= 32'h0000e2bf;
        11'h58b: sin <= 32'h0000e2d6;
        11'h58c: sin <= 32'h0000e2ee;
        11'h58d: sin <= 32'h0000e305;
        11'h58e: sin <= 32'h0000e31c;
        11'h58f: sin <= 32'h0000e333;
        11'h590: sin <= 32'h0000e34b;
        11'h591: sin <= 32'h0000e362;
        11'h592: sin <= 32'h0000e379;
        11'h593: sin <= 32'h0000e390;
        11'h594: sin <= 32'h0000e3a7;
        11'h595: sin <= 32'h0000e3be;
        11'h596: sin <= 32'h0000e3d5;
        11'h597: sin <= 32'h0000e3ec;
        11'h598: sin <= 32'h0000e403;
        11'h599: sin <= 32'h0000e419;
        11'h59a: sin <= 32'h0000e430;
        11'h59b: sin <= 32'h0000e447;
        11'h59c: sin <= 32'h0000e45e;
        11'h59d: sin <= 32'h0000e474;
        11'h59e: sin <= 32'h0000e48b;
        11'h59f: sin <= 32'h0000e4a2;
        11'h5a0: sin <= 32'h0000e4b8;
        11'h5a1: sin <= 32'h0000e4cf;
        11'h5a2: sin <= 32'h0000e4e5;
        11'h5a3: sin <= 32'h0000e4fc;
        11'h5a4: sin <= 32'h0000e512;
        11'h5a5: sin <= 32'h0000e529;
        11'h5a6: sin <= 32'h0000e53f;
        11'h5a7: sin <= 32'h0000e556;
        11'h5a8: sin <= 32'h0000e56c;
        11'h5a9: sin <= 32'h0000e582;
        11'h5aa: sin <= 32'h0000e598;
        11'h5ab: sin <= 32'h0000e5af;
        11'h5ac: sin <= 32'h0000e5c5;
        11'h5ad: sin <= 32'h0000e5db;
        11'h5ae: sin <= 32'h0000e5f1;
        11'h5af: sin <= 32'h0000e607;
        11'h5b0: sin <= 32'h0000e61d;
        11'h5b1: sin <= 32'h0000e633;
        11'h5b2: sin <= 32'h0000e649;
        11'h5b3: sin <= 32'h0000e65f;
        11'h5b4: sin <= 32'h0000e675;
        11'h5b5: sin <= 32'h0000e68b;
        11'h5b6: sin <= 32'h0000e6a1;
        11'h5b7: sin <= 32'h0000e6b7;
        11'h5b8: sin <= 32'h0000e6cc;
        11'h5b9: sin <= 32'h0000e6e2;
        11'h5ba: sin <= 32'h0000e6f8;
        11'h5bb: sin <= 32'h0000e70e;
        11'h5bc: sin <= 32'h0000e723;
        11'h5bd: sin <= 32'h0000e739;
        11'h5be: sin <= 32'h0000e74e;
        11'h5bf: sin <= 32'h0000e764;
        11'h5c0: sin <= 32'h0000e779;
        11'h5c1: sin <= 32'h0000e78f;
        11'h5c2: sin <= 32'h0000e7a4;
        11'h5c3: sin <= 32'h0000e7ba;
        11'h5c4: sin <= 32'h0000e7cf;
        11'h5c5: sin <= 32'h0000e7e4;
        11'h5c6: sin <= 32'h0000e7fa;
        11'h5c7: sin <= 32'h0000e80f;
        11'h5c8: sin <= 32'h0000e824;
        11'h5c9: sin <= 32'h0000e839;
        11'h5ca: sin <= 32'h0000e84e;
        11'h5cb: sin <= 32'h0000e864;
        11'h5cc: sin <= 32'h0000e879;
        11'h5cd: sin <= 32'h0000e88e;
        11'h5ce: sin <= 32'h0000e8a3;
        11'h5cf: sin <= 32'h0000e8b8;
        11'h5d0: sin <= 32'h0000e8cd;
        11'h5d1: sin <= 32'h0000e8e1;
        11'h5d2: sin <= 32'h0000e8f6;
        11'h5d3: sin <= 32'h0000e90b;
        11'h5d4: sin <= 32'h0000e920;
        11'h5d5: sin <= 32'h0000e935;
        11'h5d6: sin <= 32'h0000e949;
        11'h5d7: sin <= 32'h0000e95e;
        11'h5d8: sin <= 32'h0000e973;
        11'h5d9: sin <= 32'h0000e987;
        11'h5da: sin <= 32'h0000e99c;
        11'h5db: sin <= 32'h0000e9b1;
        11'h5dc: sin <= 32'h0000e9c5;
        11'h5dd: sin <= 32'h0000e9da;
        11'h5de: sin <= 32'h0000e9ee;
        11'h5df: sin <= 32'h0000ea02;
        11'h5e0: sin <= 32'h0000ea17;
        11'h5e1: sin <= 32'h0000ea2b;
        11'h5e2: sin <= 32'h0000ea3f;
        11'h5e3: sin <= 32'h0000ea54;
        11'h5e4: sin <= 32'h0000ea68;
        11'h5e5: sin <= 32'h0000ea7c;
        11'h5e6: sin <= 32'h0000ea90;
        11'h5e7: sin <= 32'h0000eaa4;
        11'h5e8: sin <= 32'h0000eab8;
        11'h5e9: sin <= 32'h0000eacc;
        11'h5ea: sin <= 32'h0000eae0;
        11'h5eb: sin <= 32'h0000eaf4;
        11'h5ec: sin <= 32'h0000eb08;
        11'h5ed: sin <= 32'h0000eb1c;
        11'h5ee: sin <= 32'h0000eb30;
        11'h5ef: sin <= 32'h0000eb44;
        11'h5f1: sin <= 32'h0000eb6c;
        11'h5f0: sin <= 32'h0000eb58;
        11'h5f3: sin <= 32'h0000eb93;
        11'h5f2: sin <= 32'h0000eb7f;
        11'h5f5: sin <= 32'h0000ebba;
        11'h5f4: sin <= 32'h0000eba7;
        11'h5f7: sin <= 32'h0000ebe2;
        11'h5f6: sin <= 32'h0000ebce;
        11'h5f9: sin <= 32'h0000ec09;
        11'h5f8: sin <= 32'h0000ebf5;
        11'h5fb: sin <= 32'h0000ec2f;
        11'h5fa: sin <= 32'h0000ec1c;
        11'h5fd: sin <= 32'h0000ec56;
        11'h5fc: sin <= 32'h0000ec43;
        11'h5ff: sin <= 32'h0000ec7d;
        11'h5fe: sin <= 32'h0000ec69;
        11'h601: sin <= 32'h0000eca3;
        11'h600: sin <= 32'h0000ec90;
        11'h603: sin <= 32'h0000ecc9;
        11'h602: sin <= 32'h0000ecb6;
        11'h605: sin <= 32'h0000ecf0;
        11'h604: sin <= 32'h0000ecdd;
        11'h607: sin <= 32'h0000ed16;
        11'h606: sin <= 32'h0000ed03;
        11'h609: sin <= 32'h0000ed3b;
        11'h608: sin <= 32'h0000ed29;
        11'h60b: sin <= 32'h0000ed61;
        11'h60a: sin <= 32'h0000ed4e;
        11'h60d: sin <= 32'h0000ed87;
        11'h60c: sin <= 32'h0000ed74;
        11'h60f: sin <= 32'h0000edac;
        11'h60e: sin <= 32'h0000ed99;
        11'h611: sin <= 32'h0000edd1;
        11'h610: sin <= 32'h0000edbf;
        11'h613: sin <= 32'h0000edf7;
        11'h612: sin <= 32'h0000ede4;
        11'h615: sin <= 32'h0000ee1c;
        11'h614: sin <= 32'h0000ee09;
        11'h617: sin <= 32'h0000ee40;
        11'h616: sin <= 32'h0000ee2e;
        11'h619: sin <= 32'h0000ee65;
        11'h618: sin <= 32'h0000ee53;
        11'h61b: sin <= 32'h0000ee8a;
        11'h61a: sin <= 32'h0000ee78;
        11'h61d: sin <= 32'h0000eeae;
        11'h61c: sin <= 32'h0000ee9c;
        11'h61f: sin <= 32'h0000eed2;
        11'h61e: sin <= 32'h0000eec0;
        11'h621: sin <= 32'h0000eef7;
        11'h620: sin <= 32'h0000eee5;
        11'h623: sin <= 32'h0000ef1b;
        11'h622: sin <= 32'h0000ef09;
        11'h625: sin <= 32'h0000ef3e;
        11'h624: sin <= 32'h0000ef2d;
        11'h627: sin <= 32'h0000ef62;
        11'h626: sin <= 32'h0000ef50;
        11'h629: sin <= 32'h0000ef86;
        11'h628: sin <= 32'h0000ef74;
        11'h62b: sin <= 32'h0000efa9;
        11'h62a: sin <= 32'h0000ef98;
        11'h62d: sin <= 32'h0000efcc;
        11'h62c: sin <= 32'h0000efbb;
        11'h62f: sin <= 32'h0000eff0;
        11'h62e: sin <= 32'h0000efde;
        11'h631: sin <= 32'h0000f013;
        11'h630: sin <= 32'h0000f001;
        11'h633: sin <= 32'h0000f035;
        11'h632: sin <= 32'h0000f024;
        11'h635: sin <= 32'h0000f058;
        11'h634: sin <= 32'h0000f047;
        11'h637: sin <= 32'h0000f07b;
        11'h636: sin <= 32'h0000f069;
        11'h639: sin <= 32'h0000f09d;
        11'h638: sin <= 32'h0000f08c;
        11'h63b: sin <= 32'h0000f0bf;
        11'h63a: sin <= 32'h0000f0ae;
        11'h63d: sin <= 32'h0000f0e1;
        11'h63c: sin <= 32'h0000f0d0;
        11'h63f: sin <= 32'h0000f103;
        11'h63e: sin <= 32'h0000f0f2;
        11'h641: sin <= 32'h0000f125;
        11'h640: sin <= 32'h0000f114;
        11'h643: sin <= 32'h0000f147;
        11'h642: sin <= 32'h0000f136;
        11'h645: sin <= 32'h0000f169;
        11'h644: sin <= 32'h0000f158;
        11'h647: sin <= 32'h0000f18a;
        11'h646: sin <= 32'h0000f179;
        11'h649: sin <= 32'h0000f1ab;
        11'h648: sin <= 32'h0000f19b;
        11'h64b: sin <= 32'h0000f1cc;
        11'h64a: sin <= 32'h0000f1bc;
        11'h64d: sin <= 32'h0000f1ed;
        11'h64c: sin <= 32'h0000f1dd;
        11'h64f: sin <= 32'h0000f20e;
        11'h64e: sin <= 32'h0000f1fe;
        11'h651: sin <= 32'h0000f22f;
        11'h650: sin <= 32'h0000f21e;
        11'h653: sin <= 32'h0000f24f;
        11'h652: sin <= 32'h0000f23f;
        11'h655: sin <= 32'h0000f270;
        11'h654: sin <= 32'h0000f25f;
        11'h657: sin <= 32'h0000f290;
        11'h656: sin <= 32'h0000f280;
        11'h659: sin <= 32'h0000f2b0;
        11'h658: sin <= 32'h0000f2a0;
        11'h65b: sin <= 32'h0000f2d0;
        11'h65a: sin <= 32'h0000f2c0;
        11'h65d: sin <= 32'h0000f2f0;
        11'h65c: sin <= 32'h0000f2e0;
        11'h65f: sin <= 32'h0000f30f;
        11'h65e: sin <= 32'h0000f2ff;
        11'h661: sin <= 32'h0000f32f;
        11'h660: sin <= 32'h0000f31f;
        11'h663: sin <= 32'h0000f34e;
        11'h662: sin <= 32'h0000f33e;
        11'h665: sin <= 32'h0000f36d;
        11'h664: sin <= 32'h0000f35e;
        11'h667: sin <= 32'h0000f38c;
        11'h666: sin <= 32'h0000f37d;
        11'h669: sin <= 32'h0000f3ab;
        11'h668: sin <= 32'h0000f39c;
        11'h66b: sin <= 32'h0000f3ca;
        11'h66a: sin <= 32'h0000f3bb;
        11'h66d: sin <= 32'h0000f3e9;
        11'h66c: sin <= 32'h0000f3d9;
        11'h66f: sin <= 32'h0000f407;
        11'h66e: sin <= 32'h0000f3f8;
        11'h671: sin <= 32'h0000f425;
        11'h670: sin <= 32'h0000f416;
        11'h673: sin <= 32'h0000f444;
        11'h672: sin <= 32'h0000f434;
        11'h675: sin <= 32'h0000f462;
        11'h674: sin <= 32'h0000f453;
        11'h677: sin <= 32'h0000f47f;
        11'h676: sin <= 32'h0000f471;
        11'h679: sin <= 32'h0000f49d;
        11'h678: sin <= 32'h0000f48e;
        11'h67b: sin <= 32'h0000f4bb;
        11'h67a: sin <= 32'h0000f4ac;
        11'h67d: sin <= 32'h0000f4d8;
        11'h67c: sin <= 32'h0000f4c9;
        11'h67f: sin <= 32'h0000f4f5;
        11'h67e: sin <= 32'h0000f4e7;
        11'h681: sin <= 32'h0000f513;
        11'h680: sin <= 32'h0000f504;
        11'h683: sin <= 32'h0000f530;
        11'h682: sin <= 32'h0000f521;
        11'h685: sin <= 32'h0000f54c;
        11'h684: sin <= 32'h0000f53e;
        11'h687: sin <= 32'h0000f569;
        11'h686: sin <= 32'h0000f55b;
        11'h689: sin <= 32'h0000f586;
        11'h688: sin <= 32'h0000f577;
        11'h68b: sin <= 32'h0000f5a2;
        11'h68a: sin <= 32'h0000f594;
        11'h68d: sin <= 32'h0000f5be;
        11'h68c: sin <= 32'h0000f5b0;
        11'h68f: sin <= 32'h0000f5da;
        11'h68e: sin <= 32'h0000f5cc;
        11'h691: sin <= 32'h0000f5f6;
        11'h690: sin <= 32'h0000f5e8;
        11'h693: sin <= 32'h0000f612;
        11'h692: sin <= 32'h0000f604;
        11'h695: sin <= 32'h0000f62e;
        11'h694: sin <= 32'h0000f620;
        11'h697: sin <= 32'h0000f649;
        11'h696: sin <= 32'h0000f63c;
        11'h699: sin <= 32'h0000f665;
        11'h698: sin <= 32'h0000f657;
        11'h69b: sin <= 32'h0000f680;
        11'h69a: sin <= 32'h0000f672;
        11'h69d: sin <= 32'h0000f69b;
        11'h69c: sin <= 32'h0000f68d;
        11'h69f: sin <= 32'h0000f6b6;
        11'h69e: sin <= 32'h0000f6a8;
        11'h6a1: sin <= 32'h0000f6d1;
        11'h6a0: sin <= 32'h0000f6c3;
        11'h6a3: sin <= 32'h0000f6eb;
        11'h6a2: sin <= 32'h0000f6de;
        11'h6a5: sin <= 32'h0000f706;
        11'h6a4: sin <= 32'h0000f6f9;
        11'h6a7: sin <= 32'h0000f720;
        11'h6a6: sin <= 32'h0000f713;
        11'h6a9: sin <= 32'h0000f73a;
        11'h6a8: sin <= 32'h0000f72d;
        11'h6ab: sin <= 32'h0000f754;
        11'h6aa: sin <= 32'h0000f747;
        11'h6ad: sin <= 32'h0000f76e;
        11'h6ac: sin <= 32'h0000f761;
        11'h6af: sin <= 32'h0000f788;
        11'h6ae: sin <= 32'h0000f77b;
        11'h6b1: sin <= 32'h0000f7a1;
        11'h6b0: sin <= 32'h0000f795;
        11'h6b3: sin <= 32'h0000f7bb;
        11'h6b2: sin <= 32'h0000f7ae;
        11'h6b5: sin <= 32'h0000f7d4;
        11'h6b4: sin <= 32'h0000f7c8;
        11'h6b7: sin <= 32'h0000f7ed;
        11'h6b6: sin <= 32'h0000f7e1;
        11'h6b9: sin <= 32'h0000f806;
        11'h6b8: sin <= 32'h0000f7fa;
        11'h6bb: sin <= 32'h0000f81f;
        11'h6ba: sin <= 32'h0000f813;
        11'h6bd: sin <= 32'h0000f838;
        11'h6bc: sin <= 32'h0000f82b;
        11'h6bf: sin <= 32'h0000f850;
        11'h6be: sin <= 32'h0000f844;
        11'h6c1: sin <= 32'h0000f869;
        11'h6c0: sin <= 32'h0000f85c;
        11'h6c3: sin <= 32'h0000f881;
        11'h6c2: sin <= 32'h0000f875;
        11'h6c5: sin <= 32'h0000f899;
        11'h6c4: sin <= 32'h0000f88d;
        11'h6c7: sin <= 32'h0000f8b1;
        11'h6c6: sin <= 32'h0000f8a5;
        11'h6c9: sin <= 32'h0000f8c9;
        11'h6c8: sin <= 32'h0000f8bd;
        11'h6cb: sin <= 32'h0000f8e0;
        11'h6ca: sin <= 32'h0000f8d4;
        11'h6cd: sin <= 32'h0000f8f8;
        11'h6cc: sin <= 32'h0000f8ec;
        11'h6cf: sin <= 32'h0000f90f;
        11'h6ce: sin <= 32'h0000f903;
        11'h6d1: sin <= 32'h0000f926;
        11'h6d0: sin <= 32'h0000f91b;
        11'h6d3: sin <= 32'h0000f93d;
        11'h6d2: sin <= 32'h0000f932;
        11'h6d5: sin <= 32'h0000f954;
        11'h6d4: sin <= 32'h0000f949;
        11'h6d7: sin <= 32'h0000f96b;
        11'h6d6: sin <= 32'h0000f960;
        11'h6d9: sin <= 32'h0000f981;
        11'h6d8: sin <= 32'h0000f976;
        11'h6db: sin <= 32'h0000f998;
        11'h6da: sin <= 32'h0000f98d;
        11'h6dd: sin <= 32'h0000f9ae;
        11'h6dc: sin <= 32'h0000f9a3;
        11'h6df: sin <= 32'h0000f9c4;
        11'h6de: sin <= 32'h0000f9b9;
        11'h6e1: sin <= 32'h0000f9da;
        11'h6e0: sin <= 32'h0000f9cf;
        11'h6e3: sin <= 32'h0000f9f0;
        11'h6e2: sin <= 32'h0000f9e5;
        11'h6e5: sin <= 32'h0000fa06;
        11'h6e4: sin <= 32'h0000f9fb;
        11'h6e7: sin <= 32'h0000fa1b;
        11'h6e6: sin <= 32'h0000fa11;
        11'h6e9: sin <= 32'h0000fa31;
        11'h6e8: sin <= 32'h0000fa26;
        11'h6eb: sin <= 32'h0000fa46;
        11'h6ea: sin <= 32'h0000fa3b;
        11'h6ed: sin <= 32'h0000fa5b;
        11'h6ec: sin <= 32'h0000fa50;
        11'h6ef: sin <= 32'h0000fa70;
        11'h6ee: sin <= 32'h0000fa65;
        11'h6f1: sin <= 32'h0000fa85;
        11'h6f0: sin <= 32'h0000fa7a;
        11'h6f3: sin <= 32'h0000fa99;
        11'h6f2: sin <= 32'h0000fa8f;
        11'h6f5: sin <= 32'h0000faae;
        11'h6f4: sin <= 32'h0000faa3;
        11'h6f7: sin <= 32'h0000fac2;
        11'h6f6: sin <= 32'h0000fab8;
        11'h6f9: sin <= 32'h0000fad6;
        11'h6f8: sin <= 32'h0000facc;
        11'h6fb: sin <= 32'h0000faea;
        11'h6fa: sin <= 32'h0000fae0;
        11'h6fd: sin <= 32'h0000fafe;
        11'h6fc: sin <= 32'h0000faf4;
        11'h6ff: sin <= 32'h0000fb12;
        11'h6fe: sin <= 32'h0000fb08;
        11'h701: sin <= 32'h0000fb25;
        11'h700: sin <= 32'h0000fb1c;
        11'h703: sin <= 32'h0000fb39;
        11'h702: sin <= 32'h0000fb2f;
        11'h705: sin <= 32'h0000fb4c;
        11'h704: sin <= 32'h0000fb42;
        11'h707: sin <= 32'h0000fb5f;
        11'h706: sin <= 32'h0000fb56;
        11'h709: sin <= 32'h0000fb72;
        11'h708: sin <= 32'h0000fb69;
        11'h70b: sin <= 32'h0000fb85;
        11'h70a: sin <= 32'h0000fb7b;
        11'h70d: sin <= 32'h0000fb97;
        11'h70c: sin <= 32'h0000fb8e;
        11'h70f: sin <= 32'h0000fbaa;
        11'h70e: sin <= 32'h0000fba1;
        11'h711: sin <= 32'h0000fbbc;
        11'h710: sin <= 32'h0000fbb3;
        11'h713: sin <= 32'h0000fbcf;
        11'h712: sin <= 32'h0000fbc5;
        11'h715: sin <= 32'h0000fbe1;
        11'h714: sin <= 32'h0000fbd8;
        11'h717: sin <= 32'h0000fbf2;
        11'h716: sin <= 32'h0000fbea;
        11'h719: sin <= 32'h0000fc04;
        11'h718: sin <= 32'h0000fbfb;
        11'h71b: sin <= 32'h0000fc16;
        11'h71a: sin <= 32'h0000fc0d;
        11'h71d: sin <= 32'h0000fc27;
        11'h71c: sin <= 32'h0000fc1e;
        11'h71f: sin <= 32'h0000fc38;
        11'h71e: sin <= 32'h0000fc30;
        11'h721: sin <= 32'h0000fc4a;
        11'h720: sin <= 32'h0000fc41;
        11'h723: sin <= 32'h0000fc5b;
        11'h722: sin <= 32'h0000fc52;
        11'h725: sin <= 32'h0000fc6b;
        11'h724: sin <= 32'h0000fc63;
        11'h727: sin <= 32'h0000fc7c;
        11'h726: sin <= 32'h0000fc74;
        11'h729: sin <= 32'h0000fc8d;
        11'h728: sin <= 32'h0000fc84;
        11'h72b: sin <= 32'h0000fc9d;
        11'h72a: sin <= 32'h0000fc95;
        11'h72d: sin <= 32'h0000fcad;
        11'h72c: sin <= 32'h0000fca5;
        11'h72f: sin <= 32'h0000fcbd;
        11'h72e: sin <= 32'h0000fcb5;
        11'h731: sin <= 32'h0000fccd;
        11'h730: sin <= 32'h0000fcc5;
        11'h733: sin <= 32'h0000fcdd;
        11'h732: sin <= 32'h0000fcd5;
        11'h735: sin <= 32'h0000fced;
        11'h734: sin <= 32'h0000fce5;
        11'h737: sin <= 32'h0000fcfc;
        11'h736: sin <= 32'h0000fcf4;
        11'h739: sin <= 32'h0000fd0b;
        11'h738: sin <= 32'h0000fd04;
        11'h73b: sin <= 32'h0000fd1a;
        11'h73a: sin <= 32'h0000fd13;
        11'h73d: sin <= 32'h0000fd29;
        11'h73c: sin <= 32'h0000fd22;
        11'h73f: sin <= 32'h0000fd38;
        11'h73e: sin <= 32'h0000fd31;
        11'h741: sin <= 32'h0000fd47;
        11'h740: sin <= 32'h0000fd40;
        11'h743: sin <= 32'h0000fd55;
        11'h742: sin <= 32'h0000fd4e;
        11'h745: sin <= 32'h0000fd64;
        11'h744: sin <= 32'h0000fd5d;
        11'h747: sin <= 32'h0000fd72;
        11'h746: sin <= 32'h0000fd6b;
        11'h749: sin <= 32'h0000fd80;
        11'h748: sin <= 32'h0000fd79;
        11'h74b: sin <= 32'h0000fd8e;
        11'h74a: sin <= 32'h0000fd87;
        11'h74d: sin <= 32'h0000fd9c;
        11'h74c: sin <= 32'h0000fd95;
        11'h74f: sin <= 32'h0000fdaa;
        11'h74e: sin <= 32'h0000fda3;
        11'h751: sin <= 32'h0000fdb7;
        11'h750: sin <= 32'h0000fdb0;
        11'h753: sin <= 32'h0000fdc4;
        11'h752: sin <= 32'h0000fdbe;
        11'h755: sin <= 32'h0000fdd1;
        11'h754: sin <= 32'h0000fdcb;
        11'h757: sin <= 32'h0000fdde;
        11'h756: sin <= 32'h0000fdd8;
        11'h759: sin <= 32'h0000fdeb;
        11'h758: sin <= 32'h0000fde5;
        11'h75b: sin <= 32'h0000fdf8;
        11'h75a: sin <= 32'h0000fdf2;
        11'h75d: sin <= 32'h0000fe05;
        11'h75c: sin <= 32'h0000fdfe;
        11'h75f: sin <= 32'h0000fe11;
        11'h75e: sin <= 32'h0000fe0b;
        11'h761: sin <= 32'h0000fe1d;
        11'h760: sin <= 32'h0000fe17;
        11'h763: sin <= 32'h0000fe29;
        11'h762: sin <= 32'h0000fe23;
        11'h765: sin <= 32'h0000fe35;
        11'h764: sin <= 32'h0000fe2f;
        11'h767: sin <= 32'h0000fe41;
        11'h766: sin <= 32'h0000fe3b;
        11'h769: sin <= 32'h0000fe4d;
        11'h768: sin <= 32'h0000fe47;
        11'h76b: sin <= 32'h0000fe58;
        11'h76a: sin <= 32'h0000fe52;
        11'h76d: sin <= 32'h0000fe63;
        11'h76c: sin <= 32'h0000fe5e;
        11'h76f: sin <= 32'h0000fe6f;
        11'h76e: sin <= 32'h0000fe69;
        11'h771: sin <= 32'h0000fe7a;
        11'h770: sin <= 32'h0000fe74;
        11'h773: sin <= 32'h0000fe85;
        11'h772: sin <= 32'h0000fe7f;
        11'h775: sin <= 32'h0000fe8f;
        11'h774: sin <= 32'h0000fe8a;
        11'h777: sin <= 32'h0000fe9a;
        11'h776: sin <= 32'h0000fe95;
        11'h779: sin <= 32'h0000fea4;
        11'h778: sin <= 32'h0000fe9f;
        11'h77b: sin <= 32'h0000feae;
        11'h77a: sin <= 32'h0000fea9;
        11'h77d: sin <= 32'h0000feb9;
        11'h77c: sin <= 32'h0000feb3;
        11'h77f: sin <= 32'h0000fec2;
        11'h77e: sin <= 32'h0000febe;
        11'h781: sin <= 32'h0000fecc;
        11'h780: sin <= 32'h0000fec7;
        11'h783: sin <= 32'h0000fed6;
        11'h782: sin <= 32'h0000fed1;
        11'h785: sin <= 32'h0000fedf;
        11'h784: sin <= 32'h0000fedb;
        11'h787: sin <= 32'h0000fee9;
        11'h786: sin <= 32'h0000fee4;
        11'h789: sin <= 32'h0000fef2;
        11'h788: sin <= 32'h0000feed;
        11'h78b: sin <= 32'h0000fefb;
        11'h78a: sin <= 32'h0000fef6;
        11'h78d: sin <= 32'h0000ff04;
        11'h78c: sin <= 32'h0000feff;
        11'h78f: sin <= 32'h0000ff0c;
        11'h78e: sin <= 32'h0000ff08;
        11'h791: sin <= 32'h0000ff15;
        11'h790: sin <= 32'h0000ff11;
        11'h793: sin <= 32'h0000ff1d;
        11'h792: sin <= 32'h0000ff19;
        11'h795: sin <= 32'h0000ff26;
        11'h794: sin <= 32'h0000ff22;
        11'h797: sin <= 32'h0000ff2e;
        11'h796: sin <= 32'h0000ff2a;
        11'h799: sin <= 32'h0000ff36;
        11'h798: sin <= 32'h0000ff32;
        11'h79b: sin <= 32'h0000ff3e;
        11'h79a: sin <= 32'h0000ff3a;
        11'h79d: sin <= 32'h0000ff45;
        11'h79c: sin <= 32'h0000ff41;
        11'h79f: sin <= 32'h0000ff4d;
        11'h79e: sin <= 32'h0000ff49;
        11'h7a1: sin <= 32'h0000ff54;
        11'h7a0: sin <= 32'h0000ff50;
        11'h7a3: sin <= 32'h0000ff5b;
        11'h7a2: sin <= 32'h0000ff58;
        11'h7a5: sin <= 32'h0000ff62;
        11'h7a4: sin <= 32'h0000ff5f;
        11'h7a7: sin <= 32'h0000ff69;
        11'h7a6: sin <= 32'h0000ff66;
        11'h7a9: sin <= 32'h0000ff70;
        11'h7a8: sin <= 32'h0000ff6c;
        11'h7ab: sin <= 32'h0000ff76;
        11'h7aa: sin <= 32'h0000ff73;
        11'h7ad: sin <= 32'h0000ff7d;
        11'h7ac: sin <= 32'h0000ff7a;
        11'h7af: sin <= 32'h0000ff83;
        11'h7ae: sin <= 32'h0000ff80;
        11'h7b1: sin <= 32'h0000ff89;
        11'h7b0: sin <= 32'h0000ff86;
        11'h7b3: sin <= 32'h0000ff8f;
        11'h7b2: sin <= 32'h0000ff8c;
        11'h7b5: sin <= 32'h0000ff95;
        11'h7b4: sin <= 32'h0000ff92;
        11'h7b7: sin <= 32'h0000ff9a;
        11'h7b6: sin <= 32'h0000ff98;
        11'h7b9: sin <= 32'h0000ffa0;
        11'h7b8: sin <= 32'h0000ff9d;
        11'h7bb: sin <= 32'h0000ffa5;
        11'h7ba: sin <= 32'h0000ffa3;
        11'h7bd: sin <= 32'h0000ffaa;
        11'h7bc: sin <= 32'h0000ffa8;
        11'h7bf: sin <= 32'h0000ffaf;
        11'h7be: sin <= 32'h0000ffad;
        11'h7c1: sin <= 32'h0000ffb4;
        11'h7c0: sin <= 32'h0000ffb2;
        11'h7c3: sin <= 32'h0000ffb9;
        11'h7c2: sin <= 32'h0000ffb7;
        11'h7c5: sin <= 32'h0000ffbe;
        11'h7c4: sin <= 32'h0000ffbb;
        11'h7c7: sin <= 32'h0000ffc2;
        11'h7c6: sin <= 32'h0000ffc0;
        11'h7c9: sin <= 32'h0000ffc6;
        11'h7c8: sin <= 32'h0000ffc4;
        11'h7cb: sin <= 32'h0000ffca;
        11'h7ca: sin <= 32'h0000ffc8;
        11'h7cd: sin <= 32'h0000ffce;
        11'h7cc: sin <= 32'h0000ffcc;
        11'h7cf: sin <= 32'h0000ffd2;
        11'h7ce: sin <= 32'h0000ffd0;
        11'h7d1: sin <= 32'h0000ffd6;
        11'h7d0: sin <= 32'h0000ffd4;
        11'h7d3: sin <= 32'h0000ffd9;
        11'h7d2: sin <= 32'h0000ffd7;
        11'h7d5: sin <= 32'h0000ffdc;
        11'h7d4: sin <= 32'h0000ffdb;
        11'h7d7: sin <= 32'h0000ffe0;
        11'h7d6: sin <= 32'h0000ffde;
        11'h7d9: sin <= 32'h0000ffe3;
        11'h7d8: sin <= 32'h0000ffe1;
        11'h7db: sin <= 32'h0000ffe5;
        11'h7da: sin <= 32'h0000ffe4;
        11'h7dd: sin <= 32'h0000ffe8;
        11'h7dc: sin <= 32'h0000ffe7;
        11'h7df: sin <= 32'h0000ffeb;
        11'h7de: sin <= 32'h0000ffe9;
        11'h7e1: sin <= 32'h0000ffed;
        11'h7e0: sin <= 32'h0000ffec;
        11'h7e3: sin <= 32'h0000ffef;
        11'h7e2: sin <= 32'h0000ffee;
        11'h7e5: sin <= 32'h0000fff1;
        11'h7e4: sin <= 32'h0000fff0;
        11'h7e7: sin <= 32'h0000fff3;
        11'h7e6: sin <= 32'h0000fff2;
        11'h7e9: sin <= 32'h0000fff5;
        11'h7e8: sin <= 32'h0000fff4;
        11'h7eb: sin <= 32'h0000fff7;
        11'h7ea: sin <= 32'h0000fff6;
        11'h7ed: sin <= 32'h0000fff8;
        11'h7ec: sin <= 32'h0000fff8;
        11'h7ef: sin <= 32'h0000fffa;
        11'h7ee: sin <= 32'h0000fff9;
        11'h7f1: sin <= 32'h0000fffb;
        11'h7f0: sin <= 32'h0000fffa;
        11'h7f3: sin <= 32'h0000fffc;
        11'h7f2: sin <= 32'h0000fffb;
        11'h7f5: sin <= 32'h0000fffd;
        11'h7f4: sin <= 32'h0000fffc;
        11'h7f7: sin <= 32'h0000fffd;
        11'h7f6: sin <= 32'h0000fffd;
        11'h7f9: sin <= 32'h0000fffe;
        11'h7f8: sin <= 32'h0000fffe;
        11'h7fb: sin <= 32'h0000fffe;
        11'h7fa: sin <= 32'h0000fffe;
        11'h7fd: sin <= 32'h0000fffe;
        11'h7fc: sin <= 32'h0000fffe;
        11'h7ff: sin <= 32'h0000fffe;
        11'h7fe: sin <= 32'h0000fffe;
      endcase
      if (signed_bit) out <= -sin;
      else out <= sin;
    end
  end
endmodule

